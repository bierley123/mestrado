TITLE UH JIRAU POWER FLOW (March/2018) 
* -------------------------------------------------------------------------------- 
* Notes: 
* TO-DO1: capacitors in shunt mode to the circuit breaker. 
* TO-DO2: ... 
* TO-DO3: ... 
* -------------------------------------------------------------------------------- 
* Models 
* A magnetic coupling 13.8kV to 525kV: 
.subckt COUPLING_525K  ( 1 3 )
*1,2: primary nodes 
*2,3: secondary nodes 
*13.8kV to 525kV 
Lsecondary ( 0 3 )  2.894612K
Lprimary ( 0 1 )  2.
K  Lsecondary  Lprimary  0.9999999
.ends COUPLING_525K
* 
*Version 3: 2 independent monophasic transformers in parallel. 
.subckt MONOPHASIC_TRANSFORMER_525K  ( 1 2 3 )
*1,0: primary A 
*2,0: primary B 
*3,0: secondary 
XTEa ( 1 3 )  COUPLING_525K
XTEb ( 2 3 )  COUPLING_525K
.ends MONOPHASIC_TRANSFORMER_525K
* 
* A magnetic coupling 13.8kV to 440V: 
.subckt MONOPHASIC_TRANSFORMER_440  ( 1 2 )
*1,0: primary nodes 
*2,0: secondary nodes 
*13.8kV to 440V 
Lsecondary ( 0 2 )  2.033186
Lprimary ( 0 1 )  2.K
K  Lsecondary  Lprimary  0.9999999
.ends MONOPHASIC_TRANSFORMER_440
* 
* A magnetic coupling where a=1: 
.subckt MONOPHASIC_REGULATOR  ( 1 2 )
*1,0: primary nodes 
*2,0: secondary nodes 
*a=1 
Lsecondary ( 0 2 )  2.K
Lprimary ( 0 1 )  2.K
K  Lsecondary  Lprimary  0.9999999
.ends MONOPHASIC_REGULATOR
* 
* LT1 and LT2: 
.subckt LT_LT1_LT2  ( 1 2 )
R_LT1_PI ( 1 2 ) COMPLEX( 1.624, 0.)
***R_LT1_PI ( 1 2 ) COMPLEX( 1.624, 28.765) 
***R_LT1_PI1 ( 1 0 ) COMPLEX( 0.,-4.05351K) 
***R_LT1_PI2 ( 2 0 ) COMPLEX( 0.,-4.05351K) 
.ends LT_LT1_LT2
* 
* 
* -------------------------------------------------------------------------------- 
* Netlist: SE MD, SE ME and SE Coletora 
R_D52A1_4 ( 170 171 )  100.n
R_D52A1_5 ( 175 176 )  100.n
R_D52A1_6 ( 166 167 )  100.n
R_D52BT_1 ( 0 0 )  1.E+12
R_D52BT_2 ( 0 0 )  1.E+12
R_D52C1_4 ( 168 163 )  100.n
R_D52C1_5 ( 173 172 )  100.n
R_D52C1_6 ( 164 162 )  100.n
R_D52G_1 ( 110 229 )  100.n
R_D52G_10 ( 115 235 )  100.n
R_D52G_11 ( 113 236 )  100.n
R_D52G_12 ( 112 237 )  100.n
R_D52G_13 ( 122 238 )  100.n
R_D52G_14 ( 121 239 )  100.n
R_D52G_15 ( 119 240 )  100.n
R_D52G_16 ( 118 241 )  100.n
R_D52G_17 ( 128 223 )  100.n
R_D52G_18 ( 127 224 )  100.n
R_D52G_19 ( 125 225 )  100.n
R_D52G_2 ( 109 228 )  100.n
R_D52G_20 ( 124 222 )  100.n
R_D52G_21 ( 200 134 )  100.n
R_D52G_22 ( 133 201 )  100.n
R_D52G_23 ( 202 131 )  100.n
R_D52G_24 ( 130 203 )  100.n
R_D52G_25 ( 140 196 )  100.n
R_D52G_26 ( 139 197 )  100.n
R_D52G_27 ( 137 198 )  100.n
R_D52G_28 ( 136 199 )  100.n
R_D52G_29 ( 221 158 )  100.n
R_D52G_3 ( 107 227 )  100.n
R_D52G_30 ( 220 157 )  100.n
R_D52G_31 ( 155 219 )  100.n
R_D52G_32 ( 218 154 )  100.n
R_D52G_33 ( 217 152 )  100.n
R_D52G_34 ( 216 151 )  100.n
R_D52G_35 ( 215 149 )  100.n
R_D52G_36 ( 214 148 )  100.n
R_D52G_37 ( 146 213 )  100.n
R_D52G_38 ( 212 145 )  100.n
R_D52G_39 ( 143 211 )  100.n
R_D52G_4 ( 106 226 )  100.n
R_D52G_40 ( 210 142 )  100.n
R_D52G_41 ( 192 98 )  100.n
R_D52G_42 ( 97 193 )  100.n
R_D52G_43 ( 194 95 )  100.n
R_D52G_44 ( 94 195 )  100.n
R_D52G_45 ( 92 209 )  100.n
R_D52G_46 ( 208 91 )  100.n
R_D52G_47 ( 89 207 )  100.n
R_D52G_48 ( 206 88 )  100.n
R_D52G_49 ( 86 205 )  100.n
R_D52G_5 ( 104 233 )  100.n
R_D52G_50 ( 84 204 )  100.n
R_D52G_6 ( 103 232 )  100.n
R_D52G_7 ( 101 231 )  100.n
R_D52G_8 ( 100 230 )  100.n
R_D52G_9 ( 116 234 )  100.n
R_D52L_1 ( 0 0 )  1.E+12
R_D52L_2 ( 0 0 )  1.E+12
R_D52L_3 ( 57 184 )  100.n
R_D52L_4 ( 0 0 )  1.E+12
R_D52L_5 ( 60 188 )  100.n
R_D52RE0_1 ( 0 0 )  1.E+12
R_D52T_1 ( 243 70 )  100.n
R_D52T_10 ( 78 252 )  100.n
R_D52T_11 ( 0 0 )  1.E+12
R_D52T_12 ( 248 159 )  100.n
R_D52T_13 ( 160 246 )  100.n
R_D52T_2 ( 245 71 )  100.n
R_D52T_3 ( 267 68 )  100.n
R_D52T_4 ( 264 67 )  100.n
R_D52T_5 ( 262 74 )  100.n
R_D52T_6 ( 75 261 )  100.n
R_D52T_7 ( 258 76 )  100.n
R_D52T_8 ( 256 80 )  100.n
R_D52T_9 ( 79 254 )  100.n
R_S57B1_1 ( 0 0 )  1.E+12
R_S57B1_2 ( 0 0 )  1.E+12
R_S57B2_1 ( 0 0 )  1.E+12
R_S57B2_2 ( 0 0 )  1.E+12
R_S57B3_1 ( 0 0 )  1.E+12
R_S57B3_2 ( 0 0 )  1.E+12
R_S57B4_1 ( 0 0 )  1.E+12
R_S57B4_2 ( 0 0 )  1.E+12
R_S57BT1_1 ( 0 0 )  1.E+12
R_S57BT1_2 ( 0 0 )  1.E+12
R_S57BT2_1 ( 0 0 )  1.E+12
R_S57BT2_2 ( 0 0 )  1.E+12
R_S57L1_1 ( 0 0 )  1.E+12
R_S57L1_2 ( 0 0 )  1.E+12
R_S57L1_3 ( 0 0 )  1.E+12
R_S57L1_4 ( 0 0 )  1.E+12
R_S57L1_5 ( 0 0 )  1.E+12
R_S57L2_1 ( 0 0 )  1.E+12
R_S57L2_2 ( 0 0 )  1.E+12
R_S57L2_3 ( 0 0 )  1.E+12
R_S57L2_4 ( 0 0 )  1.E+12
R_S57L2_5 ( 0 0 )  1.E+12
R_S57L3_1 ( 0 0 )  1.E+12
R_S57L3_2 ( 0 0 )  1.E+12
R_S57L3_3 ( 0 0 )  1.E+12
R_S57L3_4 ( 0 0 )  1.E+12
R_S57L3_5 ( 0 0 )  1.E+12
R_S57LA1_4 ( 0 0 )  1.E+12
R_S57LA1_5 ( 0 0 )  1.E+12
R_S57LA1_6 ( 0 0 )  1.E+12
R_S57T1_1 ( 0 0 )  1.E+12
R_S57T1_10 ( 0 0 )  1.E+12
R_S57T1_11 ( 0 0 )  1.E+12
R_S57T1_12 ( 0 0 )  1.E+12
R_S57T1_13 ( 0 0 )  1.E+12
R_S57T1_2 ( 0 0 )  1.E+12
R_S57T1_3 ( 0 0 )  1.E+12
R_S57T1_4 ( 0 0 )  1.E+12
R_S57T1_5 ( 0 0 )  1.E+12
R_S57T1_6 ( 0 0 )  1.E+12
R_S57T1_7 ( 0 0 )  1.E+12
R_S57T1_8 ( 0 0 )  1.E+12
R_S57T1_9 ( 0 0 )  1.E+12
R_S57T2_1 ( 0 0 )  1.E+12
R_S57T2_10 ( 0 0 )  1.E+12
R_S57T2_11 ( 0 0 )  1.E+12
R_S57T2_12 ( 0 0 )  1.E+12
R_S57T2_13 ( 0 0 )  1.E+12
R_S57T2_2 ( 0 0 )  1.E+12
R_S57T2_3 ( 0 0 )  1.E+12
R_S57T2_4 ( 0 0 )  1.E+12
R_S57T2_5 ( 0 0 )  1.E+12
R_S57T2_6 ( 0 0 )  1.E+12
R_S57T2_7 ( 0 0 )  1.E+12
R_S57T2_8 ( 0 0 )  1.E+12
R_S57T2_9 ( 0 0 )  1.E+12
R_S57T3_1 ( 0 0 )  1.E+12
R_S57T3_10 ( 0 0 )  1.E+12
R_S57T3_11 ( 0 0 )  1.E+12
R_S57T3_12 ( 0 0 )  1.E+12
R_S57T3_13 ( 0 0 )  1.E+12
R_S57T3_2 ( 0 0 )  1.E+12
R_S57T3_3 ( 0 0 )  1.E+12
R_S57T3_4 ( 0 0 )  1.E+12
R_S57T3_5 ( 0 0 )  1.E+12
R_S57T3_6 ( 0 0 )  1.E+12
R_S57T3_7 ( 0 0 )  1.E+12
R_S57T3_8 ( 0 0 )  1.E+12
R_S57T3_9 ( 0 0 )  1.E+12
R_S57TA_1 ( 0 0 )  1.E+12
R_S57TA_10 ( 0 0 )  1.E+12
R_S57TA_11 ( 0 0 )  1.E+12
R_S57TA_12 ( 0 0 )  1.E+12
R_S57TA_13 ( 0 0 )  1.E+12
R_S57TA_14 ( 0 0 )  1.E+12
R_S57TA_15 ( 0 0 )  1.E+12
R_S57TA_16 ( 0 0 )  1.E+12
R_S57TA_17 ( 0 0 )  1.E+12
R_S57TA_18 ( 0 0 )  1.E+12
R_S57TA_19 ( 0 0 )  1.E+12
R_S57TA_2 ( 0 0 )  1.E+12
R_S57TA_20 ( 0 0 )  1.E+12
R_S57TA_21 ( 0 0 )  1.E+12
R_S57TA_22 ( 0 0 )  1.E+12
R_S57TA_23 ( 0 0 )  1.E+12
R_S57TA_24 ( 0 0 )  1.E+12
R_S57TA_25 ( 0 0 )  1.E+12
R_S57TA_26 ( 0 0 )  1.E+12
R_S57TA_27 ( 0 0 )  1.E+12
R_S57TA_28 ( 0 0 )  1.E+12
R_S57TA_29 ( 0 0 )  1.E+12
R_S57TA_3 ( 0 0 )  1.E+12
R_S57TA_30 ( 0 0 )  1.E+12
R_S57TA_31 ( 0 0 )  1.E+12
R_S57TA_32 ( 0 0 )  1.E+12
R_S57TA_33 ( 0 0 )  1.E+12
R_S57TA_34 ( 0 0 )  1.E+12
R_S57TA_35 ( 0 0 )  1.E+12
R_S57TA_36 ( 0 0 )  1.E+12
R_S57TA_37 ( 0 0 )  1.E+12
R_S57TA_38 ( 0 0 )  1.E+12
R_S57TA_39 ( 0 0 )  1.E+12
R_S57TA_4 ( 0 0 )  1.E+12
R_S57TA_40 ( 0 0 )  1.E+12
R_S57TA_41 ( 0 0 )  1.E+12
R_S57TA_42 ( 0 0 )  1.E+12
R_S57TA_43 ( 0 0 )  1.E+12
R_S57TA_44 ( 0 0 )  1.E+12
R_S57TA_45 ( 0 0 )  1.E+12
R_S57TA_46 ( 0 0 )  1.E+12
R_S57TA_47 ( 0 0 )  1.E+12
R_S57TA_48 ( 0 0 )  1.E+12
R_S57TA_49 ( 0 0 )  1.E+12
R_S57TA_5 ( 0 0 )  1.E+12
R_S57TA_50 ( 0 0 )  1.E+12
R_S57TA_6 ( 0 0 )  1.E+12
R_S57TA_7 ( 0 0 )  1.E+12
R_S57TA_8 ( 0 0 )  1.E+12
R_S57TA_9 ( 0 0 )  1.E+12
R_S57TB_1 ( 0 0 )  1.E+12
R_S57TB_10 ( 0 0 )  1.E+12
R_S57TB_11 ( 0 0 )  1.E+12
R_S57TB_12 ( 0 0 )  1.E+12
R_S57TB_13 ( 0 0 )  1.E+12
R_S57TB_14 ( 0 0 )  1.E+12
R_S57TB_15 ( 0 0 )  1.E+12
R_S57TB_16 ( 0 0 )  1.E+12
R_S57TB_17 ( 0 0 )  1.E+12
R_S57TB_18 ( 0 0 )  1.E+12
R_S57TB_19 ( 0 0 )  1.E+12
R_S57TB_2 ( 0 0 )  1.E+12
R_S57TB_20 ( 0 0 )  1.E+12
R_S57TB_21 ( 0 0 )  1.E+12
R_S57TB_22 ( 0 0 )  1.E+12
R_S57TB_23 ( 0 0 )  1.E+12
R_S57TB_24 ( 0 0 )  1.E+12
R_S57TB_25 ( 0 0 )  1.E+12
R_S57TB_26 ( 0 0 )  1.E+12
R_S57TB_27 ( 0 0 )  1.E+12
R_S57TB_28 ( 0 0 )  1.E+12
R_S57TB_29 ( 0 0 )  1.E+12
R_S57TB_3 ( 0 0 )  1.E+12
R_S57TB_30 ( 0 0 )  1.E+12
R_S57TB_31 ( 0 0 )  1.E+12
R_S57TB_32 ( 0 0 )  1.E+12
R_S57TB_33 ( 0 0 )  1.E+12
R_S57TB_34 ( 0 0 )  1.E+12
R_S57TB_35 ( 0 0 )  1.E+12
R_S57TB_36 ( 0 0 )  1.E+12
R_S57TB_37 ( 0 0 )  1.E+12
R_S57TB_38 ( 0 0 )  1.E+12
R_S57TB_39 ( 0 0 )  1.E+12
R_S57TB_4 ( 0 0 )  1.E+12
R_S57TB_40 ( 0 0 )  1.E+12
R_S57TB_41 ( 0 0 )  1.E+12
R_S57TB_42 ( 0 0 )  1.E+12
R_S57TB_43 ( 0 0 )  1.E+12
R_S57TB_44 ( 0 0 )  1.E+12
R_S57TB_45 ( 0 0 )  1.E+12
R_S57TB_46 ( 0 0 )  1.E+12
R_S57TB_47 ( 0 0 )  1.E+12
R_S57TB_48 ( 0 0 )  1.E+12
R_S57TB_49 ( 0 0 )  1.E+12
R_S57TB_5 ( 0 0 )  1.E+12
R_S57TB_50 ( 0 0 )  1.E+12
R_S57TB_6 ( 0 0 )  1.E+12
R_S57TB_7 ( 0 0 )  1.E+12
R_S57TB_8 ( 0 0 )  1.E+12
R_S57TB_9 ( 0 0 )  1.E+12
R_S89A1_4 ( 171 51 )  100.n
R_S89A1_5 ( 0 0 )  1.E+12
R_S89A1_6 ( 0 0 )  1.E+12
R_S89AC1_4 ( 169 170 )  100.n
R_S89AC1_5 ( 174 175 )  100.n
R_S89AC1_6 ( 165 166 )  100.n
R_S89B1_1 ( 0 0 )  1.E+12
R_S89B1_2 ( 0 0 )  1.E+12
R_S89B2_1 ( 180 191 )  100.n
R_S89B2_2 ( 66 190 )  100.n
R_S89B3_1 ( 0 0 )  1.E+12
R_S89B3_2 ( 0 0 )  1.E+12
R_S89B4_1 ( 0 0 )  1.E+12
R_S89B4_2 ( 0 0 )  1.E+12
R_S89B5_1 ( 56 177 )  100.n
R_S89B5_2 ( 81 178 )  100.n
R_S89B6_1 ( 61 191 )  100.n
R_S89B6_2 ( 73 66 )  100.n
R_S89BTA_1 ( 179 180 )  100.n
R_S89BTA_2 ( 0 0 )  1.E+12
R_S89BTB_1 ( 65 190 )  100.n
R_S89BTB_2 ( 0 0 )  1.E+12
R_S89CA1_4 ( 168 169 )  100.n
R_S89CA1_5 ( 173 174 )  100.n
R_S89CA1_6 ( 164 165 )  100.n
R_S89CB1_4 ( 163 50 )  100.n
R_S89CB1_5 ( 50 172 )  100.n
R_S89CB1_6 ( 162 50 )  100.n
R_S89G_1 ( 229 108 )  100.n
R_S89G_10 ( 235 114 )  100.n
R_S89G_11 ( 236 111 )  100.n
R_S89G_12 ( 237 111 )  100.n
R_S89G_13 ( 238 120 )  100.n
R_S89G_14 ( 239 120 )  100.n
R_S89G_15 ( 240 117 )  100.n
R_S89G_16 ( 241 117 )  100.n
R_S89G_17 ( 223 126 )  100.n
R_S89G_18 ( 224 126 )  100.n
R_S89G_19 ( 225 123 )  100.n
R_S89G_2 ( 228 108 )  100.n
R_S89G_20 ( 222 123 )  100.n
R_S89G_21 ( 132 200 )  100.n
R_S89G_22 ( 201 132 )  100.n
R_S89G_23 ( 129 202 )  100.n
R_S89G_24 ( 129 203 )  100.n
R_S89G_25 ( 196 138 )  100.n
R_S89G_26 ( 197 138 )  100.n
R_S89G_27 ( 198 135 )  100.n
R_S89G_28 ( 199 135 )  100.n
R_S89G_29 ( 156 221 )  100.n
R_S89G_3 ( 227 105 )  100.n
R_S89G_30 ( 156 220 )  100.n
R_S89G_31 ( 219 153 )  100.n
R_S89G_32 ( 153 218 )  100.n
R_S89G_33 ( 150 217 )  100.n
R_S89G_34 ( 150 216 )  100.n
R_S89G_35 ( 147 215 )  100.n
R_S89G_36 ( 147 214 )  100.n
R_S89G_37 ( 213 144 )  100.n
R_S89G_38 ( 144 212 )  100.n
R_S89G_39 ( 211 141 )  100.n
R_S89G_4 ( 226 105 )  100.n
R_S89G_40 ( 141 210 )  100.n
R_S89G_41 ( 96 192 )  100.n
R_S89G_42 ( 193 96 )  100.n
R_S89G_43 ( 93 194 )  100.n
R_S89G_44 ( 93 195 )  100.n
R_S89G_45 ( 209 90 )  100.n
R_S89G_46 ( 90 208 )  100.n
R_S89G_47 ( 207 87 )  100.n
R_S89G_48 ( 87 206 )  100.n
R_S89G_49 ( 205 85 )  100.n
R_S89G_5 ( 233 102 )  100.n
R_S89G_50 ( 83 204 )  100.n
R_S89G_6 ( 232 102 )  100.n
R_S89G_7 ( 231 99 )  100.n
R_S89G_8 ( 230 99 )  100.n
R_S89G_9 ( 234 114 )  100.n
R_S89LA_1 ( 72 63 )  100.n
R_S89LA_2 ( 64 63 )  100.n
R_S89LA_3 ( 56 57 )  100.n
R_S89LA_4 ( 62 61 )  100.n
R_S89LA_5 ( 60 58 )  100.n
R_S89LA1_4 ( 269 169 )  100.n
R_S89LA1_5 ( 270 174 )  100.n
R_S89LA1_6 ( 268 165 )  100.n
R_S89LB_1 ( 72 69 )  100.n
R_S89LB_2 ( 0 0 )  1.E+12
R_S89LB_3 ( 178 57 )  100.n
R_S89LB_4 ( 62 73 )  100.n
R_S89LB_5 ( 60 77 )  100.n
R_S89LC_1 ( 53 186 )  100.n
R_S89LC_2 ( 0 0 )  1.E+12
R_S89LC_3 ( 52 184 )  100.n
R_S89LC_4 ( 187 189 )  100.n
R_S89LC_5 ( 3594 188 )  100.n
R_S89LE_1 ( 0 0 )  1.E+12
R_S89LE_2 ( 0 0 )  1.E+12
R_S89LE_3 ( 56 52 )  100.n
R_S89LE_4 ( 0 0 )  1.E+12
R_S89LE_5 ( 3594 58 )  100.n
R_S89RE1_4 ( 269 55 )  100.n
R_S89RE1_5 ( 270 55 )  100.n
R_S89RE1_6 ( 0 0 )  1.E+12
R_S89TA_1 ( 0 0 )  1.E+12
R_S89TA_10 ( 0 0 )  1.E+12
R_S89TA_11 ( 177 82 )  100.n
R_S89TA_12 ( 0 0 )  1.E+12
R_S89TA_13 ( 177 160 )  100.n
R_S89TA_2 ( 71 63 )  100.n
R_S89TA_3 ( 68 191 )  100.n
R_S89TA_4 ( 67 191 )  100.n
R_S89TA_5 ( 74 61 )  100.n
R_S89TA_6 ( 0 0 )  1.E+12
R_S89TA_7 ( 0 0 )  1.E+12
R_S89TA_8 ( 58 80 )  100.n
R_S89TA_9 ( 0 0 )  1.E+12
R_S89TB_1 ( 70 69 )  100.n
R_S89TB_10 ( 77 78 )  100.n
R_S89TB_11 ( 81 82 )  100.n
R_S89TB_12 ( 0 0 )  1.E+12
R_S89TB_13 ( 0 0 )  1.E+12
R_S89TB_2 ( 0 0 )  1.E+12
R_S89TB_3 ( 68 66 )  100.n
R_S89TB_4 ( 67 66 )  100.n
R_S89TB_5 ( 74 73 )  100.n
R_S89TB_6 ( 75 73 )  100.n
R_S89TB_7 ( 76 73 )  100.n
R_S89TB_8 ( 0 0 )  1.E+12
R_S89TB_9 ( 77 79 )  100.n
R_S89TC_1 ( 243 242 )  100.n
R_S89TC_10 ( 252 253 )  100.n
R_S89TC_11 ( 251 250 )  100.n
R_S89TC_12 ( 248 249 )  100.n
R_S89TC_13 ( 246 247 )  100.n
R_S89TC_2 ( 245 244 )  100.n
R_S89TC_3 ( 267 266 )  100.n
R_S89TC_4 ( 264 265 )  100.n
R_S89TC_5 ( 262 263 )  100.n
R_S89TC_6 ( 261 260 )  100.n
R_S89TC_7 ( 258 259 )  100.n
R_S89TC_8 ( 256 257 )  100.n
R_S89TC_9 ( 254 255 )  100.n
R_LT45_METER ( 3594 187 )  100.n
****** 
* Internal current source resistance: 
R_UG01 ( 0 8 )  100.n
R_UG02 ( 0 7 )  100.n
R_UG03 ( 0 9 )  100.n
R_UG04 ( 0 6 )  100.n
****** 
* Internal voltage source resistance: 
R_UG05 ( 0 4 )  100.n
R_UG06 ( 0 3 )  100.n
R_UG07 ( 0 5 )  100.n
R_UG08 ( 0 2 )  100.n
R_UG09 ( 0 12 )  100.n
R_UG10 ( 0 11 )  100.n
R_UG11 ( 0 13 )  100.n
R_UG12 ( 0 10 )  100.n
R_UG13 ( 0 16 )  100.n
R_UG14 ( 0 15 )  100.n
R_UG15 ( 0 17 )  100.n
R_UG16 ( 0 14 )  100.n
R_UG17 ( 0 20 )  100.n
R_UG18 ( 0 19 )  100.n
R_UG19 ( 0 21 )  100.n
R_UG20 ( 0 18 )  100.n
R_UG21 ( 0 24 )  100.n
R_UG22 ( 0 23 )  100.n
R_UG23 ( 0 25 )  100.n
R_UG24 ( 0 22 )  100.n
R_UG25 ( 0 28 )  100.n
R_UG26 ( 0 27 )  100.n
R_UG27 ( 0 29 )  100.n
R_UG28 ( 0 26 )  100.n
R_UG29 ( 0 32 )  100.n
R_UG30 ( 0 31 )  100.n
R_UG31 ( 0 33 )  100.n
R_UG32 ( 0 30 )  100.n
R_UG33 ( 0 36 )  100.n
R_UG34 ( 0 35 )  100.n
R_UG35 ( 0 37 )  100.n
R_UG36 ( 0 34 )  100.n
R_UG37 ( 0 40 )  100.n
R_UG38 ( 0 39 )  100.n
R_UG39 ( 0 41 )  100.n
R_UG40 ( 0 38 )  100.n
R_UG41 ( 0 44 )  100.n
R_UG42 ( 0 43 )  100.n
R_UG43 ( 0 45 )  100.n
R_UG44 ( 0 42 )  100.n
R_UG45 ( 0 48 )  100.n
R_UG46 ( 0 47 )  100.n
R_UG47 ( 0 49 )  100.n
R_UG48 ( 0 46 )  100.n
R_UG49 ( 0 161 )  100.n
R_UG50 ( 0 1 )  100.n
**** Valor da resistência no modo fonte de tensão 0.214245 
* For infinite bar load: 
****I_UG01 ( 110 8 ) COMPLEX( 1.0K, 0.) 
****I_UG02 ( 109 7 ) COMPLEX( 1.0K, 0.) 
I_UG01 ( 8 110 ) COMPLEX( 7.53066K, 7.53066K)
I_UG02 ( 7 109 ) COMPLEX( 7.53066K, 7.53066K)
I_UG03 ( 9 107 ) COMPLEX( 7.53066K, 7.53066K)
I_UG04 ( 6 106 ) COMPLEX( 7.53066K, 7.53066K)
I_UG05 ( 4 104 ) COMPLEX( 7.53066K, 0.)
I_UG06 ( 3 103 ) COMPLEX( 7.53066K, 0.)
I_UG07 ( 5 101 ) COMPLEX( 7.53066K, 0.)
I_UG08 ( 2 100 ) COMPLEX( 7.53066K, 0.)
I_UG09 ( 12 116 ) COMPLEX( 0.3623188, 0.)
I_UG10 ( 11 115 ) COMPLEX( 0.3623188, 0.)
I_UG11 ( 13 113 ) COMPLEX( 0.3623188, 0.)
I_UG12 ( 10 112 ) COMPLEX( 0.3623188, 0.)
I_UG13 ( 16 122 ) COMPLEX( 0.3623188, 0.)
I_UG14 ( 15 121 ) COMPLEX( 0.3623188, 0.)
I_UG15 ( 17 119 ) COMPLEX( 0.3623188, 0.)
I_UG16 ( 14 118 ) COMPLEX( 0.3623188, 0.)
I_UG17 ( 20 128 ) COMPLEX( 0.3623188, 0.)
I_UG18 ( 19 127 ) COMPLEX( 0.3623188, 0.)
I_UG19 ( 21 125 ) COMPLEX( 0.3623188, 0.)
I_UG20 ( 18 124 ) COMPLEX( 0.3623188, 0.)
I_UG21 ( 24 134 ) COMPLEX( 0.3623188, 0.)
I_UG22 ( 23 133 ) COMPLEX( 0.3623188, 0.)
I_UG23 ( 25 131 ) COMPLEX( 0.3623188, 0.)
I_UG24 ( 22 130 ) COMPLEX( 0.3623188, 0.)
I_UG25 ( 28 140 ) COMPLEX( 0.3623188, 0.)
I_UG26 ( 27 139 ) COMPLEX( 0.3623188, 0.)
I_UG27 ( 29 137 ) COMPLEX( 0.3623188, 0.)
I_UG28 ( 26 136 ) COMPLEX( 0.3623188, 0.)
I_UG29 ( 32 158 ) COMPLEX( 0.3623188, 0.)
I_UG30 ( 31 157 ) COMPLEX( 0.3623188, 0.)
I_UG31 ( 33 155 ) COMPLEX( 0.3623188, 0.)
I_UG32 ( 30 154 ) COMPLEX( 0.3623188, 0.)
I_UG33 ( 36 152 ) COMPLEX( 0.3623188, 0.)
I_UG34 ( 35 151 ) COMPLEX( 0.3623188, 0.)
I_UG35 ( 37 149 ) COMPLEX( 0.3623188, 0.)
I_UG36 ( 34 148 ) COMPLEX( 0.3623188, 0.)
I_UG37 ( 40 146 ) COMPLEX( 0.3623188, 0.)
I_UG38 ( 39 145 ) COMPLEX( 0.3623188, 0.)
I_UG39 ( 41 143 ) COMPLEX( 0.3623188, 0.)
I_UG40 ( 38 142 ) COMPLEX( 0.3623188, 0.)
I_UG41 ( 44 98 ) COMPLEX( 0.3623188, 0.)
I_UG42 ( 43 97 ) COMPLEX( 0.3623188, 0.)
I_UG43 ( 45 95 ) COMPLEX( 0.3623188, 0.)
I_UG44 ( 42 94 ) COMPLEX( 0.3623188, 0.)
I_UG45 ( 48 92 ) COMPLEX( 1.25511, 0.)
I_UG46 ( 47 91 ) COMPLEX( 1.25511, 0.)
I_UG47 ( 49 89 ) COMPLEX( 1.25511, 0.)
I_UG48 ( 46 88 ) COMPLEX( 10.0409K, 0.)
I_UG49 ( 161 86 ) COMPLEX( 7.53066K, 0.)
I_UG50 ( 1 84 ) COMPLEX( 7.53066K, 0.)
**** 
* For radial impedance load: 
*****V_UG05 ( 4 104 ) COMPLEX( 11.8K, 0.) 
*****V_UG06 ( 3 103 ) COMPLEX( 13.8K, 0.) 
*****V_UG07 ( 5 101 ) COMPLEX( 13.8K, 0.) 
*****V_UG08 ( 2 100 ) COMPLEX( 13.8K, 0.) 
*****V_UG09 ( 12 116 ) COMPLEX( 13.8K, 0.) 
*****V_UG10 ( 11 115 ) COMPLEX( 13.8K, 0.) 
*****V_UG11 ( 13 113 ) COMPLEX( 13.8K, 0.) 
*****V_UG12 ( 10 112 ) COMPLEX( 13.8K, 0.) 
*****V_UG13 ( 16 122 ) COMPLEX( 13.8K, 0.) 
*****V_UG14 ( 15 121 ) COMPLEX( 13.8K, 0.) 
*****V_UG15 ( 17 119 ) COMPLEX( 13.8K, 0.) 
*****V_UG16 ( 14 118 ) COMPLEX( 13.8K, 0.) 
*****V_UG17 ( 20 128 ) COMPLEX( 13.8K, 0.) 
*****V_UG18 ( 19 127 ) COMPLEX( 13.8K, 0.) 
*****V_UG19 ( 21 125 ) COMPLEX( 13.8K, 0.) 
*****V_UG20 ( 18 124 ) COMPLEX( 13.8K, 0.) 
*****V_UG21 ( 24 134 ) COMPLEX( 13.8K, 0.) 
*****V_UG22 ( 23 133 ) COMPLEX( 13.8K, 0.) 
*****V_UG23 ( 25 131 ) COMPLEX( 13.8K, 0.) 
*****V_UG24 ( 22 130 ) COMPLEX( 13.8K, 0.) 
*****V_UG25 ( 28 140 ) COMPLEX( 13.8K, 0.) 
*****V_UG26 ( 27 139 ) COMPLEX( 13.8K, 0.) 
*****V_UG27 ( 29 137 ) COMPLEX( 13.8K, 0.) 
*****V_UG28 ( 26 136 ) COMPLEX( 13.8K, 0.) 
*****V_UG29 ( 32 158 ) COMPLEX( 13.8K, 0.) 
*****V_UG30 ( 31 157 ) COMPLEX( 13.8K, 0.) 
*****V_UG31 ( 33 155 ) COMPLEX( 13.8K, 0.) 
*****V_UG32 ( 30 154 ) COMPLEX( 13.8K, 0.) 
*****V_UG33 ( 36 152 ) COMPLEX( 13.8K, 0.) 
*****V_UG34 ( 35 151 ) COMPLEX( 13.8K, 0.) 
*****V_UG35 ( 37 149 ) COMPLEX( 13.8K, 0.) 
*****V_UG36 ( 34 148 ) COMPLEX( 13.8K, 0.) 
*****V_UG37 ( 40 146 ) COMPLEX( 13.8K, 0.) 
*****V_UG38 ( 39 145 ) COMPLEX( 13.8K, 0.) 
*****V_UG39 ( 41 143 ) COMPLEX( 13.8K, 0.) 
*****V_UG40 ( 38 142 ) COMPLEX( 13.8K, 0.) 
*****V_UG41 ( 44 98 ) COMPLEX( 13.8K, 0.) 
*****V_UG42 ( 43 97 ) COMPLEX( 13.8K, 0.) 
*****V_UG43 ( 45 95 ) COMPLEX( 13.8K, 0.) 
*****V_UG44 ( 42 94 ) COMPLEX( 13.8K, 0.) 
*****V_UG45 ( 48 92 ) COMPLEX( 13.8K, 0.) 
*****V_UG46 ( 47 91 ) COMPLEX( 13.8K, 0.) 
*****V_UG47 ( 49 89 ) COMPLEX( 13.8K, 0.) 
*****V_UG48 ( 46 88 ) COMPLEX( 13.8K, 0.) 
********* Inverted phase (180.0) V_UG49 ( 161 86 ) ( 161 86 ) COMPLEX( 13.8K, 0.) 
*****V_UG49 ( 86 161 ) COMPLEX( 13.8K, 0.) 
********* Inverted phase (180.0) V_UG50 ( 1 84 ) ( 1 84 ) COMPLEX( 13.8K, 0.) 
*****V_UG50 ( 84 1 ) COMPLEX( 13.8K, 0.) 
X_T01 ( 105 108 242 )  MONOPHASIC_TRANSFORMER_525K
X_T02 ( 99 102 244 )  MONOPHASIC_TRANSFORMER_525K
X_T03 ( 111 114 266 )  MONOPHASIC_TRANSFORMER_525K
X_T04 ( 117 120 265 )  MONOPHASIC_TRANSFORMER_525K
X_T05 ( 123 126 263 )  MONOPHASIC_TRANSFORMER_525K
X_T06 ( 129 132 260 )  MONOPHASIC_TRANSFORMER_525K
X_T07 ( 135 138 259 )  MONOPHASIC_TRANSFORMER_525K
X_T08 ( 153 156 257 )  MONOPHASIC_TRANSFORMER_525K
X_T09 ( 147 150 255 )  MONOPHASIC_TRANSFORMER_525K
X_T10 ( 141 144 253 )  MONOPHASIC_TRANSFORMER_525K
X_T11 ( 93 96 250 )  MONOPHASIC_TRANSFORMER_525K
X_T12 ( 87 90 249 )  MONOPHASIC_TRANSFORMER_525K
X_T13 ( 83 85 247 )  MONOPHASIC_TRANSFORMER_525K
***R_LT3_METER ( 52 268 )  200.n 
***R_LT2_METER ( 54 270 )  200.n 
R_LT3_METER ( 3600 268 )  200.n
R_LT3_METER1 ( 52 3599 )  100.n
R_LT2_METER ( 3598 270 )  200.n
R_LT2_METER1 ( 54 3597 )  100.n
R_LT1_METER ( 3595 269 )  200.n
R_LT1_METER1 ( 53 3596 )  100.n
* 
X_LT1 ( 3596 3595 )  LT_LT1_LT2
X_LT2 ( 3597 3598 )  LT_LT1_LT2
X_LT3 ( 3599 3600 )  LT_LT1_LT2
* 
* Infinite grid/bar; power or current depend on V_Grid: 
R_Grid_SWITCH ( 50 273 )  100.n
V_Grid ( 271 0 ) COMPLEX( 302.776K,-245.06K)
* Reactance Xss at the secondary: Xss = 0.43*(525/13.8)^2 = 622.34168241966 
R_Grid ( 271 273 ) COMPLEX( 0.0144731, 622.342)
* 
* Radial. finite grid/bar: 
R_LOAD_BARRA_B ( 0 272 ) COMPLEX( 30.4697K,-217.775)
R_LOAD_BARRA_B_SWITCH ( 0 0 )  1.E+12
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA Geral 
R_S891xxQCE11 ( 274 368 )  100.n
R_S891xxQCE12 ( 275 375 )  100.n
R_D52CARGAxxQCMAC2 ( 0 353 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxQCMAC1 ( 0 525 ) COMPLEX( 387.2, 0.)
******R_D52206CARGAxxQCM10 ( 0 458 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM10 ( 0 485 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM10 ( 0 482 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM10 ( 0 483 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM10 ( 0 484 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM10 ( 0 481 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM10 ( 0 480 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM10 ( 0 478 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM10 ( 0 476 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM10 ( 0 477 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM10 ( 0 479 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM10 ( 0 475 ) COMPLEX( 387.2, 0.) 
******R_D52206CARGAxxQCM9 ( 0 421 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM9 ( 0 496 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM9 ( 0 493 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM9 ( 0 494 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM9 ( 0 495 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM9 ( 0 492 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM9 ( 0 491 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM9 ( 0 489 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM9 ( 0 487 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM9 ( 0 488 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM9 ( 0 490 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM9 ( 0 486 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM8 ( 0 612 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM8 ( 0 609 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM8 ( 0 610 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM8 ( 0 611 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM8 ( 0 608 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM8 ( 0 607 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM8 ( 0 605 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM8 ( 0 603 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM8 ( 0 604 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM8 ( 0 606 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM8 ( 0 602 ) COMPLEX( 387.2, 0.) 
******R_D52206CARGAxxQCM13 ( 0 402 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM13 ( 0 395 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM13 ( 0 406 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM13 ( 0 403 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM13 ( 0 404 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM13 ( 0 405 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM13 ( 0 401 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM13 ( 0 399 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM13 ( 0 397 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM13 ( 0 398 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM13 ( 0 400 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM13 ( 0 396 ) COMPLEX( 387.2, 0.) 
******R_D52206CARGAxxQCM12 ( 0 407 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM12 ( 0 418 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM12 ( 0 415 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM12 ( 0 416 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM12 ( 0 417 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM12 ( 0 414 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM12 ( 0 413 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM12 ( 0 411 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM12 ( 0 409 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM12 ( 0 410 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM12 ( 0 412 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM12 ( 0 408 ) COMPLEX( 387.2, 0.) 
******R_D52205CARGAxxQCM11 ( 0 543 ) COMPLEX( 387.2, 0.) 
******R_D52204CARGAxxQCM11 ( 0 540 ) COMPLEX( 387.2, 0.) 
******R_D52203CARGAxxQCM11 ( 0 541 ) COMPLEX( 387.2, 0.) 
******R_D52202CARGAxxQCM11 ( 0 542 ) COMPLEX( 387.2, 0.) 
******R_D52201CARGAxxQCM11 ( 0 539 ) COMPLEX( 387.2, 0.) 
******R_D52106CARGAxxQCM11 ( 0 538 ) COMPLEX( 387.2, 0.) 
******R_D52105CARGAxxQCM11 ( 0 536 ) COMPLEX( 387.2, 0.) 
******R_D52104CARGAxxQCM11 ( 0 534 ) COMPLEX( 387.2, 0.) 
******R_D52103CARGAxxQCM11 ( 0 535 ) COMPLEX( 387.2, 0.) 
******R_D52102CARGAxxQCM11 ( 0 537 ) COMPLEX( 387.2, 0.) 
******R_D52101CARGAxxQCM11 ( 0 533 ) COMPLEX( 387.2, 0.) 
R_D52CARGAxxTSVT2 ( 0 320 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxCDTSB4 ( 0 276 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxTSVT1 ( 0 342 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxCDTSB3 ( 0 277 ) COMPLEX( 387.2, 0.)
*******R_D52206CARGAxxQCM7 ( 0 544 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM7 ( 0 554 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM7 ( 0 552 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM7 ( 0 553 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM7 ( 0 551 ) COMPLEX( 387.2, 0.) 
*******R_D52106CARGAxxQCM7 ( 0 550 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM7 ( 0 548 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM7 ( 0 546 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM7 ( 0 547 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM7 ( 0 549 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM7 ( 0 545 ) COMPLEX( 387.2, 0.) 
*******R_D52206CARGAxxQCM6 ( 0 555 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM6 ( 0 566 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM6 ( 0 563 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM6 ( 0 564 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM6 ( 0 565 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM6 ( 0 562 ) COMPLEX( 387.2, 0.) 
*******R_D52106CARGAxxQCM6 ( 0 561 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM6 ( 0 559 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM6 ( 0 557 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM6 ( 0 558 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM6 ( 0 560 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM6 ( 0 556 ) COMPLEX( 387.2, 0.) 
*******R_D52206CARGAxxQCM5 ( 0 567 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM5 ( 0 578 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM5 ( 0 575 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM5 ( 0 576 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM5 ( 0 577 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM5 ( 0 574 ) COMPLEX( 387.2, 0.) 
*******R_D52106CARGAxxQCM5 ( 0 573 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM5 ( 0 571 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM5 ( 0 569 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM5 ( 0 570 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM5 ( 0 572 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM5 ( 0 568 ) COMPLEX( 387.2, 0.) 
R_D52CARGAxxQCME2 ( 0 432 ) COMPLEX( 387.2, 0.)
*******R_D52205CARGAxxQCM4 ( 0 622 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM4 ( 0 619 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM4 ( 0 620 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM4 ( 0 621 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM4 ( 0 618 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM4 ( 0 616 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM4 ( 0 614 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM4 ( 0 615 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM4 ( 0 617 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM4 ( 0 613 ) COMPLEX( 387.2, 0.) 
*******R_D52206CARGAxxQCM3 ( 0 590 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM3 ( 0 601 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM3 ( 0 598 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM3 ( 0 599 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM3 ( 0 600 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM3 ( 0 597 ) COMPLEX( 387.2, 0.) 
*******R_D52106CARGAxxQCM3 ( 0 596 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM3 ( 0 594 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM3 ( 0 592 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM3 ( 0 593 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM3 ( 0 595 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM3 ( 0 591 ) COMPLEX( 387.2, 0.) 
*******R_D52206CARGAxxQCM2 ( 0 454 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM2 ( 0 589 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM2 ( 0 586 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM2 ( 0 587 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM2 ( 0 588 ) COMPLEX( 387.2, 0.) 
*******R_D52201CARGAxxQCM2 ( 0 585 ) COMPLEX( 387.2, 0.) 
*******R_D52106CARGAxxQCM2 ( 0 584 ) COMPLEX( 387.2, 0.) 
*******R_D52105CARGAxxQCM2 ( 0 582 ) COMPLEX( 387.2, 0.) 
*******R_D52104CARGAxxQCM2 ( 0 580 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM2 ( 0 581 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM2 ( 0 583 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM2 ( 0 579 ) COMPLEX( 387.2, 0.) 
*******R_D52205CARGAxxQCM1 ( 0 638 ) COMPLEX( 387.2, 0.) 
*******R_D52204CARGAxxQCM1 ( 0 635 ) COMPLEX( 387.2, 0.) 
*******R_D52203CARGAxxQCM1 ( 0 636 ) COMPLEX( 387.2, 0.) 
*******R_D52202CARGAxxQCM1 ( 0 637 ) COMPLEX( 387.2, 0.) 
***********R_D52106CARGAxxQCM1 ( 0 633 ) COMPLEX( 387.2, 0.) 
*******R_D52103CARGAxxQCM1 ( 0 629 ) COMPLEX( 387.2, 0.) 
*******R_D52102CARGAxxQCM1 ( 0 632 ) COMPLEX( 387.2, 0.) 
*******R_D52101CARGAxxQCM1 ( 0 625 ) COMPLEX( 387.2, 0.) 
R_D52QLxxQCM11 ( 364 365 )  100.n
X_TSE3 ( 516 511 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM8 ( 443 444 )  100.n
X_TSB2 ( 456 529 )  MONOPHASIC_REGULATOR
X_TSE2 ( 522 526 )  MONOPHASIC_TRANSFORMER_440
R_D52QEExxQCM2 ( 526 455 )  100.n
R_D52QE1xxQCM2 ( 531 455 )  100.n
X_TSA3 ( 530 531 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM2 ( 455 453 )  100.n
R_D52QE2xxQCM2 ( 532 453 )  100.n
X_TSA4 ( 528 532 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM1 ( 623 624 )  100.n
R_D52xxQCGE1 ( 0 0 )  1.E+12
R_D52xxQCGE2 ( 0 0 )  1.E+12
R_D52xxCDG26 ( 0 0 )  1.E+12
R_D52xxCDG25 ( 85 386 )  100.n
X_TSA26 ( 387 388 )  MONOPHASIC_TRANSFORMER_440
X_TSA25 ( 386 385 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM13 ( 388 389 )  100.n
R_D52QE1xxQCM13 ( 385 390 )  100.n
R_D52QEExxQCM13 ( 384 390 )  100.n
R_D52QLxxQCM13 ( 389 390 )  100.n
X_TSE13 ( 383 384 )  MONOPHASIC_TRANSFORMER_440
R_S891xxQCE13 ( 382 383 )  100.n
R_S892xxQCE13 ( 374 382 )  100.n
R_S893xxQCE13 ( 0 0 )  1.E+12
R_D52206xxQCM13 ( 389 402 )  100.n
R_D52204xxQCM13 ( 389 406 )  100.n
R_D52205xxQCM13 ( 395 389 )  100.n
R_D52203xxQCM13 ( 389 403 )  100.n
R_D52202xxQCM13 ( 389 404 )  100.n
R_D52201xxQCM13 ( 405 389 )  100.n
R_D52106xxQCM13 ( 390 401 )  100.n
R_D52105xxQCM13 ( 390 399 )  100.n
R_D52104xxQCM13 ( 390 397 )  100.n
R_D52103xxQCM13 ( 0 0 )  1.E+12
R_D52102xxQCM13 ( 390 400 )  100.n
R_D52101xxQCM13 ( 396 390 )  100.n
R_D52QLxxQCM12 ( 362 363 )  100.n
X_TSE7 ( 335 327 )  MONOPHASIC_TRANSFORMER_440
X_TSB4 ( 322 323 )  MONOPHASIC_REGULATOR
R_D52xxCDTSB4 ( 0 0 )  1.E+12
R_D52ExxCDG14E ( 135 324 )  100.n
R_D522xxCDG14S ( 0 0 )  1.E+12
R_D521xxCDG14S ( 0 0 )  1.E+12
R_D52xxCDG13 ( 138 326 )  100.n
R_D52QLxxQCM7 ( 331 330 )  100.n
X_TSA14 ( 325 328 )  MONOPHASIC_TRANSFORMER_440
X_TSA13 ( 326 329 )  MONOPHASIC_TRANSFORMER_440
X_TSVT2 ( 320 321 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM7 ( 328 330 )  100.n
R_D52QE1xxQCM7 ( 329 331 )  100.n
R_D52QEExxQCM7 ( 327 331 )  100.n
R_D52206xxQCM7 ( 0 0 )  1.E+12
R_D52204xxQCM7 ( 0 0 )  1.E+12
R_D52205xxQCM7 ( 330 554 )  100.n
R_D52203xxQCM7 ( 552 330 )  100.n
R_D52202xxQCM7 ( 330 553 )  100.n
R_D52201xxQCM7 ( 330 551 )  100.n
R_D52106xxQCM7 ( 331 550 )  100.n
R_D52105xxQCM7 ( 331 548 )  100.n
R_D52104xxQCM7 ( 331 546 )  100.n
R_D52103xxQCM7 ( 547 331 )  100.n
R_D52102xxQCM7 ( 331 549 )  100.n
R_D52101xxQCM7 ( 0 0 )  1.E+12
R_D52207xxQCM6 ( 0 0 )  1.E+12
X_TSVT1 ( 342 341 )  MONOPHASIC_TRANSFORMER_440
X_TSE6 ( 337 338 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDTSB3 ( 0 0 )  1.E+12
X_TSB3 ( 348 349 )  MONOPHASIC_REGULATOR
R_D522xxCDG12S ( 347 348 )  100.n
R_D521xxCDG12S ( 346 347 )  100.n
R_D52ExxCDG12E ( 0 0 )  1.E+12
X_TSA12 ( 346 345 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM6 ( 345 343 )  100.n
R_D52QE1xxQCM6 ( 340 344 )  100.n
R_D52QEExxQCM6 ( 338 344 )  100.n
R_D52QLxxQCM6 ( 344 343 )  100.n
X_TSA11 ( 339 340 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG11 ( 132 339 )  100.n
R_D52206xxQCM6 ( 343 555 )  100.n
R_D52204xxQCM6 ( 0 0 )  1.E+12
R_D52205xxQCM6 ( 343 566 )  100.n
R_D52203xxQCM6 ( 564 343 )  100.n
R_D52202xxQCM6 ( 343 565 )  100.n
R_D52201xxQCM6 ( 343 562 )  100.n
R_D52106xxQCM6 ( 344 561 )  100.n
R_D52105xxQCM6 ( 344 559 )  100.n
R_D52104xxQCM6 ( 344 557 )  100.n
R_D52103xxQCM6 ( 558 344 )  100.n
R_D52102xxQCM6 ( 344 560 )  100.n
R_D52101xxQCM6 ( 0 0 )  1.E+12
R_D52206xxQCM5 ( 449 567 )  100.n
R_D52205xxQCM5 ( 449 578 )  100.n
R_D52201xxQCM5 ( 449 574 )  100.n
R_D52204xxQCM5 ( 0 0 )  1.E+12
R_D52203xxQCM5 ( 576 449 )  100.n
R_D52202xxQCM5 ( 449 577 )  100.n
R_D52106xxQCM5 ( 450 573 )  100.n
R_D52QLxxQCM5 ( 450 449 )  100.n
R_D52105xxQCM5 ( 450 571 )  100.n
R_D52104xxQCM5 ( 450 569 )  100.n
R_D52103xxQCM5 ( 570 450 )  100.n
R_D52102xxQCM5 ( 450 572 )  100.n
R_D52101xxQCM5 ( 0 0 )  1.E+12
X_TSE5 ( 333 315 )  MONOPHASIC_TRANSFORMER_440
* X_TSG1 ( 351 437 ) MONOPHASIC_TRANSFORMER_440 
X_TSG1 ( 437 351 )  MONOPHASIC_TRANSFORMER_440
X_TSG2 ( 436 350 )  MONOPHASIC_TRANSFORMER_440
R_S892xxQCE11 ( 366 274 )  100.n
R_S893xxQCE11 ( 0 0 )  1.E+12
X_TSE11 ( 368 369 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM11 ( 373 364 )  100.n
R_D52QEExxQCM11 ( 369 365 )  100.n
R_D52QE1xxQCM11 ( 370 365 )  100.n
X_TSA21 ( 371 370 )  MONOPHASIC_TRANSFORMER_440
X_TSA22 ( 372 373 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG21 ( 96 371 )  100.n
R_D52xxCDG22 ( 0 0 )  1.E+12
V_UGD7 ( 391 0 ) COMPLEX( 440., 0.)
R_D52xxQCGE7 ( 0 0 )  1.E+12
X_TSG7 ( 393 392 )  MONOPHASIC_TRANSFORMER_440
R_D522xxQCME4 ( 393 394 )  100.n
R_D523xxQCME4 ( 394 381 )  100.n
R_D521xxQCME4 ( 394 439 )  100.n
R_D52QLxxQCM3 ( 425 424 )  100.n
R_D52QEExxQCM3 ( 511 425 )  100.n
R_D52QE1xxQCM3 ( 513 425 )  100.n
X_TSA5 ( 521 513 )  MONOPHASIC_TRANSFORMER_440
X_TSA6 ( 514 512 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM3 ( 512 424 )  100.n
R_D52QEExxQCM4 ( 504 452 )  100.n
R_D52QE1xxQCM4 ( 506 452 )  100.n
X_TSE4 ( 509 504 )  MONOPHASIC_TRANSFORMER_440
X_TSA7 ( 510 506 )  MONOPHASIC_TRANSFORMER_440
X_TSB6 ( 441 459 )  MONOPHASIC_REGULATOR
R_D52QLxxQCM10 ( 419 420 )  100.n
R_D52QLxxQCM9 ( 422 423 )  100.n
R_D52QLxxQCM4 ( 452 451 )  100.n
R_D52QE2xxQCM4 ( 505 451 )  100.n
X_TSA8 ( 507 505 )  MONOPHASIC_TRANSFORMER_440
R_S891xxQCE8 ( 502 503 )  100.n
R_S892xxQCE8 ( 440 502 )  100.n
R_S893xxQCE8 ( 0 0 )  1.E+12
R_D52106xxQCM11 ( 365 538 )  100.n
R_D52104xxQCM11 ( 365 534 )  100.n
R_D52105xxQCM11 ( 365 536 )  100.n
R_D52201xxQCM11 ( 364 539 )  100.n
R_D52202xxQCM11 ( 542 364 )  100.n
R_D52203xxQCM11 ( 364 541 )  100.n
R_D52204xxQCM11 ( 364 540 )  100.n
R_D52205xxQCM11 ( 364 543 )  100.n
R_D52103xxQCM11 ( 0 0 )  1.E+12
R_D52102xxQCM11 ( 365 537 )  100.n
R_D52101xxQCM11 ( 533 365 )  100.n
R_D52106xxQCM12 ( 363 413 )  100.n
R_D52104xxQCM12 ( 363 409 )  100.n
R_D52105xxQCM12 ( 363 411 )  100.n
R_D52201xxQCM12 ( 362 414 )  100.n
R_D52202xxQCM12 ( 417 362 )  100.n
R_D52203xxQCM12 ( 362 416 )  100.n
R_D52204xxQCM12 ( 362 415 )  100.n
R_D52205xxQCM12 ( 362 418 )  100.n
R_D52206xxQCM12 ( 407 362 )  100.n
R_D52103xxQCM12 ( 0 0 )  1.E+12
R_D52102xxQCM12 ( 363 412 )  100.n
R_D52101xxQCM12 ( 408 363 )  100.n
R_S893xxQCE12 ( 0 0 )  1.E+12
R_S892xxQCE12 ( 367 275 )  100.n
X_TSE12 ( 375 376 )  MONOPHASIC_TRANSFORMER_440
R_D52QEExxQCM12 ( 376 363 )  100.n
R_D52QE1xxQCM12 ( 377 363 )  100.n
R_D52QE2xxQCM12 ( 380 362 )  100.n
X_TSA24 ( 379 380 )  MONOPHASIC_TRANSFORMER_440
X_TSA23 ( 378 377 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG24 ( 0 0 )  1.E+12
R_D52xxCDG23 ( 90 378 )  100.n
V_UGD5 ( 355 0 ) COMPLEX( 440., 0.)
V_UGD6 ( 356 0 ) COMPLEX( 440., 0.)
R_D52xxQCGE5 ( 0 0 )  1.E+12
R_D52xxQCGE6 ( 0 0 )  1.E+12
X_TSG5 ( 360 357 )  MONOPHASIC_TRANSFORMER_440
X_TSG6 ( 359 358 )  MONOPHASIC_TRANSFORMER_440
R_D525xxQCME3 ( 361 439 )  100.n
R_D522xxQCME3 ( 361 440 )  100.n
R_D524xxQCME3 ( 359 361 )  100.n
R_D523xxQCME3 ( 360 361 )  100.n
R_D521xxQCME3 ( 0 0 )  1.E+12
R_D525Q1xxQCMAC2 ( 353 441 )  100.n
R_D524Q1xxQCMAC2 ( 353 354 )  100.n
R_D522Q1xxQCMAC2 ( 354 445 )  100.n
R_D525xxQCME2 ( 307 435 )  100.n
R_D521xxQCME2 ( 435 427 )  100.n
R_D524xxQCME2 ( 432 435 )  100.n
R_D523xxQCME2 ( 0 0 )  1.E+12
R_D522xxQCME2 ( 0 0 )  1.E+12
X_TSG3 ( 434 430 )  MONOPHASIC_TRANSFORMER_440
X_TSG4 ( 433 431 )  MONOPHASIC_TRANSFORMER_440
R_D52xxQCGE3 ( 0 0 )  1.E+12
R_D52xxQCGE4 ( 0 0 )  1.E+12
V_UGD4 ( 428 0 ) COMPLEX( 440., 0.)
V_UGD3 ( 429 0 ) COMPLEX( 440., 0.)
V_UGD2 ( 352 0 ) COMPLEX( 440., 0.)
V_UGD1 ( 527 0 ) COMPLEX( 440., 0.)
R_D524xxQCME1 ( 0 0 )  1.E+12
R_D523xxQCME1 ( 0 0 )  1.E+12
R_D525xxQCME1 ( 427 438 )  100.n
R_D522xxQCME1 ( 0 0 )  1.E+12
R_D521xxQCME1 ( 0 0 )  1.E+12
R_D524Q1xxQCMAC1 ( 314 525 )  100.n
R_D525Q1xxQCMAC1 ( 525 456 )  100.n
R_D522Q1xxQCMAC1 ( 524 314 )  100.n
R_D52ExxCDG20E ( 0 0 )  1.E+12
R_D522xxCDG20S ( 0 0 )  1.E+12
R_D521xxCDG20S ( 460 461 )  100.n
R_D52xxCDG19 ( 144 467 )  100.n
X_TSA20 ( 461 463 )  MONOPHASIC_TRANSFORMER_440
X_TSA19 ( 467 464 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM10 ( 463 419 )  100.n
R_D52QE1xxQCM10 ( 464 420 )  100.n
R_D52QEExxQCM10 ( 462 420 )  100.n
R_D52206xxQCM10 ( 419 458 )  100.n
R_D52204xxQCM10 ( 419 482 )  100.n
R_D52205xxQCM10 ( 0 0 )  1.E+12
R_D52203xxQCM10 ( 419 483 )  100.n
R_D52202xxQCM10 ( 484 419 )  100.n
R_D52201xxQCM10 ( 419 481 )  100.n
R_D52106xxQCM10 ( 420 480 )  100.n
R_D52105xxQCM10 ( 420 478 )  100.n
R_D52104xxQCM10 ( 420 476 )  100.n
R_D52103xxQCM10 ( 477 420 )  100.n
R_D52102xxQCM10 ( 420 479 )  100.n
R_D52101xxQCM10 ( 475 420 )  100.n
R_D52xxCDG18 ( 0 0 )  1.E+12
R_D52xxCDG17 ( 150 474 )  100.n
R_S892xxQCE9 ( 442 472 )  100.n
R_S893xxQCE9 ( 0 0 )  1.E+12
R_S891xxQCE9 ( 472 473 )  100.n
R_S892xxQCE10 ( 457 465 )  100.n
R_S893xxQCE10 ( 0 0 )  1.E+12
R_S891xxQCE10 ( 465 466 )  100.n
X_TSE10 ( 466 462 )  MONOPHASIC_TRANSFORMER_440
X_TSE9 ( 473 468 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM9 ( 469 422 )  100.n
X_TSA18 ( 471 469 )  MONOPHASIC_TRANSFORMER_440
X_TSA17 ( 474 470 )  MONOPHASIC_TRANSFORMER_440
R_D52QE1xxQCM9 ( 470 423 )  100.n
R_D52QEExxQCM9 ( 468 423 )  100.n
R_D52206xxQCM9 ( 421 422 )  100.n
R_D52204xxQCM9 ( 422 493 )  100.n
R_D52205xxQCM9 ( 422 496 )  100.n
R_D52203xxQCM9 ( 422 494 )  100.n
R_D52202xxQCM9 ( 495 422 )  100.n
R_D52201xxQCM9 ( 422 492 )  100.n
R_D52106xxQCM9 ( 423 491 )  100.n
R_D52105xxQCM9 ( 423 489 )  100.n
R_D52104xxQCM9 ( 423 487 )  100.n
R_D52103xxQCM9 ( 488 423 )  100.n
R_D52102xxQCM9 ( 423 490 )  100.n
R_D52101xxQCM9 ( 486 423 )  100.n
X_TSB5 ( 445 447 )  MONOPHASIC_REGULATOR
X_TSE8 ( 503 497 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM8 ( 498 443 )  100.n
R_D52QE1xxQCM8 ( 499 444 )  100.n
R_D52QEExxQCM8 ( 497 444 )  100.n
X_TSA16 ( 500 498 )  MONOPHASIC_TRANSFORMER_440
X_TSA15 ( 448 499 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG16 ( 0 0 )  1.E+12
R_D522xxCDG15S ( 446 448 )  100.n
R_D521xxCDG15S ( 0 0 )  1.E+12
R_D52ExxCDG15E ( 156 446 )  100.n
R_D52xxCDG8 ( 0 0 )  1.E+12
R_D52xxCDG7 ( 120 510 )  100.n
R_D52xxCDG6 ( 0 0 )  1.E+12
R_D52xxCDG5 ( 114 521 )  100.n
R_D52206xxQCM2 ( 454 453 )  100.n
R_D52204xxQCM2 ( 0 0 )  1.E+12
R_D52205xxQCM2 ( 453 589 )  100.n
R_D52203xxQCM2 ( 587 453 )  100.n
R_D52202xxQCM2 ( 453 588 )  100.n
R_D52201xxQCM2 ( 453 585 )  100.n
R_D52106xxQCM2 ( 455 584 )  100.n
R_D52105xxQCM2 ( 455 582 )  100.n
R_D52104xxQCM2 ( 455 580 )  100.n
R_D52103xxQCM2 ( 581 455 )  100.n
R_D52102xxQCM2 ( 455 583 )  100.n
R_D52101xxQCM2 ( 579 455 )  100.n
R_D52QE2xxQCM5 ( 318 449 )  100.n
R_D52QE1xxQCM5 ( 319 450 )  100.n
R_D52QEExxQCM5 ( 315 450 )  100.n
X_TSA10 ( 317 318 )  MONOPHASIC_TRANSFORMER_440
X_TSA9 ( 316 319 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG10 ( 0 0 )  1.E+12
R_D52xxCDG9 ( 126 316 )  100.n
R_S893xxQCE6 ( 0 0 )  1.E+12
R_C574xxQCE6 ( 0 0 )  1.E+12
R_S892xxQCE6 ( 0 0 )  1.E+12
R_C573xxQCE6 ( 0 0 )  1.E+12
R_C572xxQCE6 ( 0 0 )  1.E+12
R_S891xxQCE6 ( 336 337 )  100.n
R_C571xxQCE6 ( 0 0 )  1.E+12
R_S893xxQCE7 ( 0 0 )  1.E+12
R_C574xxQCE7 ( 0 0 )  1.E+12
R_S892xxQCE7 ( 307 334 )  100.n
R_C573xxQCE7 ( 0 0 )  1.E+12
R_C572xxQCE7 ( 0 0 )  1.E+12
R_S891xxQCE7 ( 334 335 )  100.n
R_C571xxQCE7 ( 0 0 )  1.E+12
R_S893xxQCE5 ( 0 0 )  1.E+12
R_C574xxQCE5 ( 0 0 )  1.E+12
R_S892xxQCE5 ( 0 0 )  1.E+12
R_C573xxQCE5 ( 0 0 )  1.E+12
R_C572xxQCE5 ( 0 0 )  1.E+12
R_S891xxQCE5 ( 332 333 )  100.n
R_C571xxQCE5 ( 0 0 )  1.E+12
R_S893xxQCE2 ( 0 0 )  1.E+12
R_C574xxQCE2 ( 0 0 )  1.E+12
R_S892xxQCE2 ( 0 0 )  1.E+12
R_C573xxQCE2 ( 0 0 )  1.E+12
R_C572xxQCE2 ( 0 0 )  1.E+12
R_S891xxQCE2 ( 520 522 )  100.n
R_C571xxQCE2 ( 0 0 )  1.E+12
R_S893xxQCE3 ( 0 0 )  1.E+12
R_C574xxQCE3 ( 0 0 )  1.E+12
R_S892xxQCE3 ( 0 0 )  1.E+12
R_C573xxQCE3 ( 0 0 )  1.E+12
R_C572xxQCE3 ( 0 0 )  1.E+12
R_S891xxQCE3 ( 515 516 )  100.n
R_C571xxQCE3 ( 0 0 )  1.E+12
R_S893xxQCE4 ( 0 0 )  1.E+12
R_C574xxQCE4 ( 0 0 )  1.E+12
R_S892xxQCE4 ( 0 0 )  1.E+12
R_C573xxQCE4 ( 0 0 )  1.E+12
R_C572xxQCE4 ( 0 0 )  1.E+12
R_S891xxQCE4 ( 508 509 )  100.n
R_C571xxQCE4 ( 0 0 )  1.E+12
R_S893xxQCE1 ( 312 517 )  100.n
R_C574xxQCE1 ( 0 0 )  1.E+12
R_S892xxQCE1 ( 0 0 )  1.E+12
R_C573xxQCE1 ( 0 0 )  1.E+12
R_C572xxQCE1 ( 0 0 )  1.E+12
R_S891xxQCE1 ( 517 518 )  100.n
R_C571xxQCE1 ( 0 0 )  1.E+12
X_TSE1 ( 518 519 )  MONOPHASIC_TRANSFORMER_440
R_D52201xxQCM3 ( 424 597 )  100.n
R_D52205xxQCM3 ( 424 601 )  100.n
R_D52206xxQCM3 ( 0 0 )  1.E+12
R_D52204xxQCM3 ( 424 598 )  100.n
R_D52203xxQCM3 ( 599 424 )  100.n
R_D52202xxQCM3 ( 424 600 )  100.n
R_D52106xxQCM3 ( 425 596 )  100.n
R_D52105xxQCM3 ( 425 594 )  100.n
R_D52104xxQCM3 ( 425 592 )  100.n
R_D52103xxQCM3 ( 593 425 )  100.n
R_D52102xxQCM3 ( 425 595 )  100.n
R_D52101xxQCM3 ( 0 0 )  1.E+12
R_D52204xxQCM4 ( 0 0 )  1.E+12
R_D52205xxQCM4 ( 451 622 )  100.n
R_D52203xxQCM4 ( 620 451 )  100.n
R_D52202xxQCM4 ( 451 621 )  100.n
R_D52201xxQCM4 ( 451 618 )  100.n
R_D52105xxQCM4 ( 452 616 )  100.n
R_D52104xxQCM4 ( 452 614 )  100.n
R_D52103xxQCM4 ( 615 452 )  100.n
R_D52102xxQCM4 ( 452 617 )  100.n
R_D52101xxQCM4 ( 0 0 )  1.E+12
R_D52204xxQCM8 ( 443 609 )  100.n
R_D52205xxQCM8 ( 443 612 )  100.n
R_D52203xxQCM8 ( 443 610 )  100.n
R_D52202xxQCM8 ( 611 443 )  100.n
R_D52201xxQCM8 ( 443 608 )  100.n
R_D52106xxQCM8 ( 444 607 )  100.n
R_D52105xxQCM8 ( 444 605 )  100.n
R_D52104xxQCM8 ( 444 603 )  100.n
R_D52103xxQCM8 ( 604 444 )  100.n
R_D52102xxQCM8 ( 444 606 )  100.n
R_D52101xxQCM8 ( 602 444 )  100.n
R_D52204xxQCM1 ( 0 0 )  1.E+12
R_D52205xxQCM1 ( 624 638 )  100.n
R_D52203xxQCM1 ( 624 636 )  100.n
R_D52202xxQCM1 ( 637 624 )  100.n
R_D52201xxQCM1 ( 624 634 )  100.n
R_D52106xxQCM1 ( 623 633 )  100.n
R_D52105xxQCM1 ( 623 630 )  100.n
R_D52104xxQCM1 ( 623 626 )  100.n
R_D52103xxQCM1 ( 629 623 )  100.n
R_D52102xxQCM1 ( 623 632 )  100.n
R_D52101xxQCM1 ( 0 0 )  1.E+12
R_D52QEExxQCM1 ( 519 623 )  100.n
R_D52QE2xxQCM1 ( 631 624 )  100.n
R_D52QE1xxQCM1 ( 628 623 )  100.n
X_TSA2 ( 627 631 )  MONOPHASIC_TRANSFORMER_440
X_TSA1 ( 523 628 )  MONOPHASIC_TRANSFORMER_440
X_TSB1 ( 426 524 )  MONOPHASIC_REGULATOR
R_D52ExxCDG3E ( 102 302 )  100.n
R_D522xxCDG3S ( 302 530 )  100.n
R_D521xxCDG3S ( 0 0 )  1.E+12
R_D52xxCDG4 ( 0 0 )  1.E+12
R_D52xxCDG2 ( 0 0 )  1.E+12
R_D521xxCDG1S ( 0 0 )  1.E+12
R_D522xxCDG1S ( 303 523 )  100.n
R_D52ExxCDG1E ( 108 303 )  100.n
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG1 
R_D52322LOADxxQSG1 ( 639 0 ) COMPLEX( 59.048, 0.)
R_D52322xxQSG1 ( 639 640 )  100.n
R_D52323LOADxxQSG1 ( 641 0 ) COMPLEX( 2.4495,-0.8052)
R_D52323xxQSG1 ( 641 640 )  100.n
R_D52321LOADxxQSG1 ( 0 642 ) COMPLEX( 20.4906,-13.2357)
R_D52321xxQSG1 ( 642 640 )  100.n
R_D52320LOADxxQSG1 ( 0 643 ) COMPLEX( 20.4906,-13.2357)
R_D52320xxQSG1 ( 640 643 )  100.n
R_D52307xxQSG1 ( 644 640 )  100.n
R_D52307LOADxxQSG1 ( 644 0 ) COMPLEX( 390., 0.)
R_D52309xxQSG1 ( 645 640 )  100.n
R_D52309LOADxxQSG1 ( 0 645 ) COMPLEX( 390., 0.)
R_D52319LOADxxQSG1 ( 646 0 ) COMPLEX( 390., 0.)
R_D52319xxQSG1 ( 646 640 )  100.n
R_D52318LOADxxQSG1 ( 647 0 ) COMPLEX( 6.078,-3.2805)
R_D52318xxQSG1 ( 647 640 )  100.n
R_D52310LOADxxQSG1 ( 648 0 ) COMPLEX( 390., 0.)
R_D52310xxQSG1 ( 648 640 )  100.n
R_D52317LOADxxQSG1 ( 649 0 ) COMPLEX( 6.078,-3.2805)
R_D52317xxQSG1 ( 649 640 )  100.n
R_D52316LOADxxQSG1 ( 650 0 ) COMPLEX( 123.9039,-92.928)
R_D52316xxQSG1 ( 650 640 )  100.n
R_D52315LOADxxQSG1 ( 651 0 ) COMPLEX( 2.4495,-0.8052)
R_D52315xxQSG1 ( 651 640 )  100.n
R_D52314LOADxxQSG1 ( 652 0 ) COMPLEX( 390., 0.)
R_D52314xxQSG1 ( 652 640 )  100.n
R_D52313LOADxxQSG1 ( 653 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG1 ( 653 640 )  100.n
R_D52312LOADxxQSG1 ( 654 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG1 ( 654 640 )  100.n
R_D52311LOADxxQSG1 ( 655 0 ) COMPLEX( 20.4906,-13.2357)
R_D52311xxQSG1 ( 655 640 )  100.n
R_D52308xxQSG1 ( 656 640 )  100.n
R_D52308LOADxxQSG1 ( 0 656 ) COMPLEX( 59.048, 0.)
R_D52306LOADxxQSG1 ( 0 657 ) COMPLEX( 2.4495,-0.8052)
R_D52306xxQSG1 ( 657 640 )  100.n
R_D52305LOADxxQSG1 ( 0 658 ) COMPLEX( 59.048, 0.)
R_D52305xxQSG1 ( 658 640 )  100.n
R_D52304LOADxxQSG1 ( 0 659 ) COMPLEX( 390., 0.)
R_D52304xxQSG1 ( 659 640 )  100.n
R_D52303LOADxxQSG1 ( 0 660 ) COMPLEX( 176.6793,-141.7467)
R_D52303xxQSG1 ( 660 640 )  100.n
R_D52302LOADxxQSG1 ( 0 661 ) COMPLEX( 390., 0.)
R_D52302xxQSG1 ( 661 640 )  100.n
R_D52301LOADxxQSG1 ( 0 662 ) COMPLEX( 2.0445,-1.1034)
R_D52301xxQSG1 ( 640 662 )  100.n
R_D52207xxQSG1 ( 664 665 )  100.n
R_D52207LOADxxQSG1 ( 664 0 ) COMPLEX( 390., 0.)
R_D52209xxQSG1 ( 666 665 )  100.n
R_D52209LOADxxQSG1 ( 0 666 ) COMPLEX( 4.773,-2.832)
R_D52219LOADxxQSG1 ( 667 0 ) COMPLEX( 3.9963,-2.265)
R_D52219xxQSG1 ( 667 665 )  100.n
R_D52218LOADxxQSG1 ( 668 0 ) COMPLEX( 3.9963,-2.265)
R_D52218xxQSG1 ( 668 665 )  100.n
R_D52210LOADxxQSG1 ( 669 0 ) COMPLEX( 390., 0.)
R_D52210xxQSG1 ( 669 665 )  100.n
R_D52217LOADxxQSG1 ( 670 0 ) COMPLEX( 390., 0.)
R_D52217xxQSG1 ( 670 665 )  100.n
R_D52216LOADxxQSG1 ( 671 0 ) COMPLEX( 390., 0.)
R_D52216xxQSG1 ( 671 665 )  100.n
R_D52215LOADxxQSG1 ( 672 0 ) COMPLEX( 13.9875,-8.6688)
R_D52215xxQSG1 ( 672 665 )  100.n
R_D52214LOADxxQSG1 ( 673 0 ) COMPLEX( 16.3926,-10.5885)
R_D52214xxQSG1 ( 673 665 )  100.n
R_D52213LOADxxQSG1 ( 674 0 ) COMPLEX( 235.5726,-188.9955)
R_D52213xxQSG1 ( 674 665 )  100.n
R_D52212LOADxxQSG1 ( 675 0 ) COMPLEX( 38.148,-23.6421)
R_D52212xxQSG1 ( 675 665 )  100.n
R_D52211LOADxxQSG1 ( 676 0 ) COMPLEX( 390., 0.)
R_D52211xxQSG1 ( 676 665 )  100.n
R_D52208xxQSG1 ( 677 665 )  100.n
R_D52208LOADxxQSG1 ( 0 677 ) COMPLEX( 59.048, 0.)
R_D52206LOADxxQSG1 ( 663 678 )  100.n
R_D52206xxQSG1 ( 678 665 )  100.n
R_D52205LOADxxQSG1 ( 0 679 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG1 ( 679 665 )  100.n
R_D52204LOADxxQSG1 ( 0 680 ) COMPLEX( 3.9963,-2.265)
R_D52204xxQSG1 ( 680 665 )  100.n
R_D52203LOADxxQSG1 ( 0 681 ) COMPLEX( 123.9039,-92.928)
R_D52203xxQSG1 ( 681 665 )  100.n
R_D52202LOADxxQSG1 ( 0 682 ) COMPLEX( 86.7843,-60.576)
R_D52202xxQSG1 ( 682 665 )  100.n
R_D52201LOADxxQSG1 ( 0 683 ) COMPLEX( 38.148,-23.6421)
R_D52201xxQSG1 ( 665 683 )  100.n
R_D52E1xxQSG1 ( 626 687 )  100.n
R_D52E2xxQSG1 ( 585 665 )  100.n
R_D52L2xxQSG1 ( 640 665 )  100.n
R_D52107xxQSG1 ( 686 687 )  100.n
R_D52107LOADxxQSG1 ( 0 0 )  1.E+12
R_D52109xxQSG1 ( 688 687 )  100.n
R_D52109LOADxxQSG1 ( 0 688 ) COMPLEX( 3.9963,-2.265)
R_D52119LOADxxQSG1 ( 689 0 ) COMPLEX( 3.9963,-2.265)
R_D52119xxQSG1 ( 689 687 )  100.n
R_D52118LOADxxQSG1 ( 690 0 ) COMPLEX( 16.3926,-10.5885)
R_D52118xxQSG1 ( 690 687 )  100.n
R_D52110LOADxxQSG1 ( 691 0 ) COMPLEX( 16.3926,-10.5885)
R_D52110xxQSG1 ( 691 687 )  100.n
R_D52117LOADxxQSG1 ( 692 0 ) COMPLEX( 390., 0.)
R_D52117xxQSG1 ( 692 687 )  100.n
R_D52L1xxQSG1 ( 0 0 )  1.E+12
R_D52116LOADxxQSG1 ( 694 0 ) COMPLEX( 13.9875,-8.6688)
R_D52116xxQSG1 ( 694 687 )  100.n
R_D52115LOADxxQSG1 ( 695 0 ) COMPLEX( 235.5726,-188.9955)
R_D52115xxQSG1 ( 695 687 )  100.n
R_D52114LOADxxQSG1 ( 696 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG1 ( 696 687 )  100.n
R_D52113LOADxxQSG1 ( 697 0 ) COMPLEX( 4.773,-2.832)
R_D52113xxQSG1 ( 697 687 )  100.n
R_D52112LOADxxQSG1 ( 698 0 ) COMPLEX( 53.3484,-35.8503)
R_D52112xxQSG1 ( 698 687 )  100.n
R_D52111LOADxxQSG1 ( 699 0 ) COMPLEX( 390., 0.)
R_D52111xxQSG1 ( 699 687 )  100.n
R_D52108xxQSG1 ( 700 687 )  100.n
R_D52108LOADxxQSG1 ( 0 700 ) COMPLEX( 390., 0.)
R_D52106LOADxxQSG1 ( 0 701 ) COMPLEX( 20.4906,-13.2357)
R_D52106xxQSG1 ( 701 687 )  100.n
R_D52105LOADxxQSG1 ( 0 702 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG1 ( 702 687 )  100.n
R_D52104LOADxxQSG1 ( 0 703 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG1 ( 703 687 )  100.n
R_D52103LOADxxQSG1 ( 0 704 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG1 ( 704 687 )  100.n
R_D52102LOADxxQSG1 ( 0 705 ) COMPLEX( 390., 0.)
R_D52102xxQSG1 ( 705 687 )  100.n
R_D52101LOADxxQSG1 ( 0 706 ) COMPLEX( 53.3484,-35.8503)
R_D52101xxQSG1 ( 687 706 )  100.n
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG2 
R_D52207xxQSG2 ( 708 709 )  100.n
R_D52207LOADxxQSG2 ( 708 0 ) COMPLEX( 390., 0.)
R_D52209xxQSG2 ( 710 709 )  100.n
R_D52209LOADxxQSG2 ( 0 710 ) COMPLEX( 390., 0.)
R_D52210LOADxxQSG2 ( 711 0 ) COMPLEX( 390., 0.)
R_D52210xxQSG2 ( 711 709 )  100.n
R_D52216LOADxxQSG2 ( 712 0 ) COMPLEX( 3.9963,-2.265)
R_D52216xxQSG2 ( 712 709 )  100.n
R_D52215LOADxxQSG2 ( 713 0 ) COMPLEX( 390., 0.)
R_D52215xxQSG2 ( 713 709 )  100.n
R_D52214LOADxxQSG2 ( 714 0 ) COMPLEX( 16.3926,-10.5885)
R_D52214xxQSG2 ( 714 709 )  100.n
R_D52213LOADxxQSG2 ( 715 0 ) COMPLEX( 235.5726,-188.9955)
R_D52213xxQSG2 ( 715 709 )  100.n
R_D52212LOADxxQSG2 ( 716 0 ) COMPLEX( 390., 0.)
R_D52212xxQSG2 ( 716 709 )  100.n
R_D52211LOADxxQSG2 ( 717 0 ) COMPLEX( 49.368, 0.)
R_D52211xxQSG2 ( 717 709 )  100.n
R_D52208xxQSG2 ( 718 709 )  100.n
R_D52208LOADxxQSG2 ( 0 718 ) COMPLEX( 390., 0.)
R_D52206LOADxxQSG2 ( 707 719 )  100.n
R_D52206xxQSG2 ( 719 709 )  100.n
R_D52205LOADxxQSG2 ( 0 720 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG2 ( 720 709 )  100.n
R_D52204LOADxxQSG2 ( 0 721 ) COMPLEX( 3.9963,-2.265)
R_D52204xxQSG2 ( 721 709 )  100.n
R_D52203LOADxxQSG2 ( 0 722 ) COMPLEX( 123.9039,-92.928)
R_D52203xxQSG2 ( 722 709 )  100.n
R_D52202LOADxxQSG2 ( 0 723 ) COMPLEX( 86.7843,-60.576)
R_D52202xxQSG2 ( 723 709 )  100.n
R_D52201LOADxxQSG2 ( 0 724 ) COMPLEX( 49.368, 0.)
R_D52201xxQSG2 ( 709 724 )  100.n
R_D52307xxQSG2 ( 725 726 )  100.n
R_D52307LOADxxQSG2 ( 725 0 ) COMPLEX( 2.4495,-0.8052)
R_D52309xxQSG2 ( 727 726 )  100.n
R_D52309LOADxxQSG2 ( 0 727 ) COMPLEX( 390., 0.)
R_D52319LOADxxQSG2 ( 728 0 ) COMPLEX( 390., 0.)
R_D52319xxQSG2 ( 728 726 )  100.n
R_D52318LOADxxQSG2 ( 729 0 ) COMPLEX( 20.4906,-13.2357)
R_D52318xxQSG2 ( 729 726 )  100.n
R_D52310LOADxxQSG2 ( 730 0 ) COMPLEX( 168.96,-126.72)
R_D52310xxQSG2 ( 730 726 )  100.n
R_D52317LOADxxQSG2 ( 731 0 ) COMPLEX( 20.4906,-13.2357)
R_D52317xxQSG2 ( 731 726 )  100.n
R_D52316LOADxxQSG2 ( 732 0 ) COMPLEX( 6.078,-3.2805)
R_D52316xxQSG2 ( 732 726 )  100.n
R_D52315LOADxxQSG2 ( 733 0 ) COMPLEX( 390., 0.)
R_D52315xxQSG2 ( 733 726 )  100.n
R_D52314LOADxxQSG2 ( 734 0 ) COMPLEX( 6.078,-3.2805)
R_D52314xxQSG2 ( 734 726 )  100.n
R_D52313LOADxxQSG2 ( 735 0 ) COMPLEX( 390., 0.)
R_D52313xxQSG2 ( 735 726 )  100.n
R_D52312LOADxxQSG2 ( 736 0 ) COMPLEX( 64.2471,-51.5442)
R_D52312xxQSG2 ( 736 726 )  100.n
R_D52311LOADxxQSG2 ( 737 0 ) COMPLEX( 390., 0.)
R_D52311xxQSG2 ( 737 726 )  100.n
R_D52308xxQSG2 ( 738 726 )  100.n
R_D52308LOADxxQSG2 ( 0 738 ) COMPLEX( 20.4906,-13.2357)
R_D52306LOADxxQSG2 ( 0 739 ) COMPLEX( 2.4495,-0.8052)
R_D52306xxQSG2 ( 739 726 )  100.n
R_D52305LOADxxQSG2 ( 0 740 ) COMPLEX( 390., 0.)
R_D52305xxQSG2 ( 740 726 )  100.n
R_D52304LOADxxQSG2 ( 0 741 ) COMPLEX( 20.4906,-13.2357)
R_D52304xxQSG2 ( 741 726 )  100.n
R_D52303LOADxxQSG2 ( 0 742 ) COMPLEX( 6.078,-3.2805)
R_D52303xxQSG2 ( 742 726 )  100.n
R_D52302LOADxxQSG2 ( 0 743 ) COMPLEX( 390., 0.)
R_D52302xxQSG2 ( 743 726 )  100.n
R_D52301LOADxxQSG2 ( 0 744 ) COMPLEX( 2.0445,-1.1034)
R_D52301xxQSG2 ( 726 744 )  100.n
R_D52E1xxQSG2 ( 580 748 )  100.n
R_D52E2xxQSG2 ( 634 709 )  100.n
R_D52L2xxQSG2 ( 726 709 )  100.n
R_D52107xxQSG2 ( 747 748 )  100.n
R_D52107LOADxxQSG2 ( 747 0 ) COMPLEX( 390., 0.)
R_D52109xxQSG2 ( 749 748 )  100.n
R_D52109LOADxxQSG2 ( 0 749 ) COMPLEX( 3.9963,-2.265)
R_D52110LOADxxQSG2 ( 750 0 ) COMPLEX( 235.5726,-188.9955)
R_D52110xxQSG2 ( 750 748 )  100.n
R_D52L1xxQSG2 ( 0 0 )  1.E+12
R_D52116LOADxxQSG2 ( 752 0 ) COMPLEX( 3.9963,-2.265)
R_D52116xxQSG2 ( 752 748 )  100.n
R_D52115LOADxxQSG2 ( 753 0 ) COMPLEX( 3.9963,-2.265)
R_D52115xxQSG2 ( 753 748 )  100.n
R_D52114LOADxxQSG2 ( 754 0 ) COMPLEX( 49.368, 0.)
R_D52114xxQSG2 ( 754 748 )  100.n
R_D52113LOADxxQSG2 ( 755 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG2 ( 755 748 )  100.n
R_D52112LOADxxQSG2 ( 756 0 ) COMPLEX( 390., 0.)
R_D52112xxQSG2 ( 756 748 )  100.n
R_D52111LOADxxQSG2 ( 757 0 ) COMPLEX( 16.3926,-10.5885)
R_D52111xxQSG2 ( 0 0 )  1.E+12
R_D52108xxQSG2 ( 758 748 )  100.n
R_D52108LOADxxQSG2 ( 0 758 ) COMPLEX( 3.9963,-2.265)
R_D52106LOADxxQSG2 ( 746 759 )  100.n
R_D52106xxQSG2 ( 759 748 )  100.n
R_D52105LOADxxQSG2 ( 0 760 ) COMPLEX( 390., 0.)
R_D52105xxQSG2 ( 760 748 )  100.n
R_D52104LOADxxQSG2 ( 0 761 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG2 ( 761 748 )  100.n
R_D52103LOADxxQSG2 ( 0 762 ) COMPLEX( 3.9963,-2.265)
R_D52103xxQSG2 ( 762 748 )  100.n
R_D52102LOADxxQSG2 ( 0 763 ) COMPLEX( 86.7843,-60.576)
R_D52102xxQSG2 ( 763 748 )  100.n
R_D52101LOADxxQSG2 ( 0 764 ) COMPLEX( 390., 0.)
R_D52101xxQSG2 ( 748 764 )  100.n
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U01CCM 
R_D52132LOADxxU01 ( 765 0 ) COMPLEX( 390., 0.)
R_D52132xxU01 ( 0 0 )  1.E+12
R_D52131LOADxxU01 ( 767 0 ) COMPLEX( 220.8492,-177.1833)
R_D52131xxU01 ( 767 766 )  100.n
R_D52130LOADxxU01 ( 769 0 ) COMPLEX( 390., 0.)
R_D52130xxU01 ( 0 0 )  1.E+12
R_D52129LOADxxU01 ( 770 0 ) COMPLEX( 390., 0.)
R_D52129xxU01 ( 0 0 )  1.E+12
R_D52128LOADxxU01 ( 771 0 ) COMPLEX( 390., 0.)
R_D52128xxU01 ( 0 0 )  1.E+12
R_D52127LOADxxU01 ( 772 0 ) COMPLEX( 76.5744,-53.4492)
R_D52127xxU01 ( 772 766 )  100.n
R_D52126LOADxxU01 ( 773 0 ) COMPLEX( 390., 0.)
R_D52126xxU01 ( 0 0 )  1.E+12
R_D52125LOADxxU01 ( 774 0 ) COMPLEX( 390., 0.)
R_D52125xxU01 ( 0 0 )  1.E+12
R_D52124xxU01 ( 775 766 )  100.n
R_D52117xxU01 ( 776 766 )  100.n
R_D52117LOADxxU01 ( 0 776 ) COMPLEX( 1.363267K,-1.593835K)
R_D52124LOADxxU01 ( 0 775 ) COMPLEX( 176.6793,-141.7467)
R_D52123LOADxxU01 ( 0 777 ) COMPLEX( 390., 0.)
R_D52123xxU01 ( 0 0 )  1.E+12
R_D52122LOADxxU01 ( 0 778 ) COMPLEX( 390., 0.)
R_D52122xxU01 ( 0 0 )  1.E+12
R_D52121LOADxxU01 ( 0 779 ) COMPLEX( 95.2656,-68.9712)
R_D52121xxU01 ( 779 766 )  100.n
R_D52120LOADxxU01 ( 0 780 ) COMPLEX( 390., 0.)
R_D52120xxU01 ( 0 0 )  1.E+12
R_D52119LOADxxU01 ( 0 781 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU01 ( 781 766 )  100.n
R_D52118LOADxxU01 ( 0 783 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU01 ( 766 783 )  100.n
R_D52115LOADxxU01 ( 784 0 ) COMPLEX( 69.7374,-48.6771)
R_D52115xxU01 ( 784 766 )  100.n
R_D52ExxU01 ( 630 766 )  100.n
R_D52116LOADxxU01 ( 786 0 ) COMPLEX( 390., 0.)
R_D52116xxU01 ( 0 0 )  1.E+12
R_D52114LOADxxU01 ( 787 0 ) COMPLEX( 69.7374,-48.6771)
R_D52114xxU01 ( 787 766 )  100.n
R_D52113LOADxxU01 ( 788 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU01 ( 788 766 )  100.n
R_D52112LOADxxU01 ( 789 0 ) COMPLEX( 3.9963,-2.265)
R_D52112xxU01 ( 789 766 )  100.n
R_D52111LOADxxU01 ( 790 0 ) COMPLEX( 390., 0.)
R_D52111xxU01 ( 0 0 )  1.E+12
R_D52110LOADxxU01 ( 791 0 ) COMPLEX( 8.1777,-4.4139)
R_D52110xxU01 ( 791 766 )  100.n
R_D52109LOADxxU01 ( 792 0 ) COMPLEX( 390., 0.)
R_D52109xxU01 ( 0 0 )  1.E+12
R_D52107xxU01 ( 793 766 )  100.n
R_D52108xxU01 ( 794 766 )  100.n
R_D52108LOADxxU01 ( 0 794 ) COMPLEX( 13.9875,-8.6688)
R_D52107LOADxxU01 ( 0 793 ) COMPLEX( 13.9875,-8.6688)
R_D52106LOADxxU01 ( 0 795 ) COMPLEX( 390., 0.)
R_D52106xxU01 ( 0 0 )  1.E+12
R_D52105LOADxxU01 ( 0 796 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU01 ( 796 766 )  100.n
R_D52104LOADxxU01 ( 0 797 ) COMPLEX( 26.6742,-17.9253)
R_D52104xxU01 ( 797 766 )  100.n
R_D52103LOADxxU01 ( 0 798 ) COMPLEX( 390., 0.)
R_D52103xxU01 ( 0 0 )  1.E+12
R_D52102LOADxxU01 ( 0 799 ) COMPLEX( 390., 0.)
R_D52102xxU01 ( 0 0 )  1.E+12
R_D52101LOADxxU01 ( 0 800 ) COMPLEX( 2.8263,-1.8255)
R_D52101xxU01 ( 766 800 )  100.n
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U02CCM 
R_D52132LOADxxU02 ( 801 0 ) COMPLEX( 390., 0.)
R_D52132xxU02 ( 0 0 )  1.E+12
R_D52131LOADxxU02 ( 803 0 ) COMPLEX( 220.8492,-177.1833)
R_D52131xxU02 ( 803 802 )  100.n
R_D52130LOADxxU02 ( 804 0 ) COMPLEX( 390., 0.)
R_D52130xxU02 ( 0 0 )  1.E+12
R_D52129LOADxxU02 ( 805 0 ) COMPLEX( 390., 0.)
R_D52129xxU02 ( 0 0 )  1.E+12
R_D52128LOADxxU02 ( 806 0 ) COMPLEX( 390., 0.)
R_D52128xxU02 ( 0 0 )  1.E+12
R_D52127LOADxxU02 ( 807 0 ) COMPLEX( 76.5744,-53.4492)
R_D52127xxU02 ( 807 802 )  100.n
R_D52126LOADxxU02 ( 808 0 ) COMPLEX( 390., 0.)
R_D52126xxU02 ( 0 0 )  1.E+12
R_D52125LOADxxU02 ( 809 0 ) COMPLEX( 390., 0.)
R_D52125xxU02 ( 0 0 )  1.E+12
R_D52124xxU02 ( 810 802 )  100.n
R_D52117xxU02 ( 811 802 )  100.n
R_D52117LOADxxU02 ( 0 811 ) COMPLEX( 1.363267K,-1.593835K)
R_D52124LOADxxU02 ( 0 810 ) COMPLEX( 176.6793,-141.7467)
R_D52123LOADxxU02 ( 0 812 ) COMPLEX( 390., 0.)
R_D52123xxU02 ( 0 0 )  1.E+12
R_D52122LOADxxU02 ( 0 813 ) COMPLEX( 390., 0.)
R_D52122xxU02 ( 0 0 )  1.E+12
R_D52121LOADxxU02 ( 0 814 ) COMPLEX( 95.2656,-68.9712)
R_D52121xxU02 ( 814 802 )  100.n
R_D52120LOADxxU02 ( 0 815 ) COMPLEX( 390., 0.)
R_D52120xxU02 ( 0 0 )  1.E+12
R_D52119LOADxxU02 ( 0 816 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU02 ( 816 802 )  100.n
R_D52118LOADxxU02 ( 0 817 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU02 ( 802 817 )  100.n
R_D52115LOADxxU02 ( 818 0 ) COMPLEX( 69.7374,-48.6771)
R_D52115xxU02 ( 818 802 )  100.n
R_D52ExxU02 ( 633 802 )  100.n
R_D52116LOADxxU02 ( 820 0 ) COMPLEX( 390., 0.)
R_D52116xxU02 ( 0 0 )  1.E+12
R_D52114LOADxxU02 ( 821 0 ) COMPLEX( 69.7374,-48.6771)
R_D52114xxU02 ( 821 802 )  100.n
R_D52113LOADxxU02 ( 822 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU02 ( 822 802 )  100.n
R_D52112LOADxxU02 ( 823 0 ) COMPLEX( 3.9963,-2.265)
R_D52112xxU02 ( 823 802 )  100.n
R_D52111LOADxxU02 ( 824 0 ) COMPLEX( 390., 0.)
R_D52111xxU02 ( 0 0 )  1.E+12
R_D52110LOADxxU02 ( 825 0 ) COMPLEX( 8.1777,-4.4139)
R_D52110xxU02 ( 825 802 )  100.n
R_D52109LOADxxU02 ( 826 0 ) COMPLEX( 390., 0.)
R_D52109xxU02 ( 0 0 )  1.E+12
R_D52107xxU02 ( 827 802 )  100.n
R_D52108xxU02 ( 828 802 )  100.n
R_D52108LOADxxU02 ( 0 828 ) COMPLEX( 13.9875,-8.6688)
R_D52107LOADxxU02 ( 0 827 ) COMPLEX( 13.9875,-8.6688)
R_D52106LOADxxU02 ( 0 829 ) COMPLEX( 390., 0.)
R_D52106xxU02 ( 0 0 )  1.E+12
R_D52105LOADxxU02 ( 0 830 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU02 ( 830 802 )  100.n
R_D52104LOADxxU02 ( 0 831 ) COMPLEX( 26.6742,-17.9253)
R_D52104xxU02 ( 831 802 )  100.n
R_D52103LOADxxU02 ( 0 832 ) COMPLEX( 390., 0.)
R_D52103xxU02 ( 0 0 )  1.E+12
R_D52102LOADxxU02 ( 0 833 ) COMPLEX( 390., 0.)
R_D52102xxU02 ( 0 0 )  1.E+12
R_D52101LOADxxU02 ( 0 834 ) COMPLEX( 2.8263,-1.8255)
R_D52101xxU02 ( 802 834 )  100.n
*------------------------------------------------------------------------------------------------------------------------ 
* Netlist: Auxiliares CA U03CCM 
R_D52132LOADxxU03 ( 835 0 ) COMPLEX( 390., 0.)
R_D52132xxU03 ( 835 836 )  1.E+12
R_D52131LOADxxU03 ( 837 0 ) COMPLEX( 220.8492,-177.1833)
R_D52131xxU03 ( 837 836 )  100.n
R_D52130LOADxxU03 ( 838 0 ) COMPLEX( 390., 0.)
R_D52130xxU03 ( 838 836 )  1.E+12
R_D52129LOADxxU03 ( 839 0 ) COMPLEX( 390., 0.)
R_D52129xxU03 ( 839 836 )  1.E+12
R_D52128LOADxxU03 ( 840 0 ) COMPLEX( 390., 0.)
R_D52128xxU03 ( 840 836 )  1.E+12
R_D52127LOADxxU03 ( 841 0 ) COMPLEX( 76.5744,-53.4492)
R_D52127xxU03 ( 841 836 )  100.n
R_D52126LOADxxU03 ( 842 0 ) COMPLEX( 390., 0.)
R_D52126xxU03 ( 842 836 )  1.E+12
R_D52125LOADxxU03 ( 843 0 ) COMPLEX( 390., 0.)
R_D52125xxU03 ( 843 836 )  1.E+12
R_D52124xxU03 ( 844 836 )  100.n
R_D52117xxU03 ( 845 836 )  100.n
R_D52117LOADxxU03 ( 0 845 ) COMPLEX( 1.363267K,-1.593835K)
R_D52124LOADxxU03 ( 0 844 ) COMPLEX( 176.6793,-141.7467)
R_D52123LOADxxU03 ( 0 846 ) COMPLEX( 390., 0.)
R_D52123xxU03 ( 846 836 )  1.E+12
R_D52122LOADxxU03 ( 0 847 ) COMPLEX( 390., 0.)
R_D52122xxU03 ( 847 836 )  1.E+12
R_D52121LOADxxU03 ( 0 848 ) COMPLEX( 95.2656,-68.9712)
R_D52121xxU03 ( 848 836 )  100.n
R_D52120LOADxxU03 ( 0 849 ) COMPLEX( 390., 0.)
R_D52120xxU03 ( 849 836 )  1.E+12
R_D52119LOADxxU03 ( 0 850 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU03 ( 850 836 )  100.n
R_D52118LOADxxU03 ( 0 851 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU03 ( 836 851 )  100.n
R_D52115LOADxxU03 ( 852 0 ) COMPLEX( 69.7374,-48.6771)
R_D52115xxU03 ( 852 836 )  100.n
R_D52ExxU03 ( 637 836 )  100.n
R_D52116LOADxxU03 ( 854 0 ) COMPLEX( 390., 0.)
R_D52116xxU03 ( 854 836 )  1.E+12
R_D52114LOADxxU03 ( 855 0 ) COMPLEX( 69.7374,-48.6771)
R_D52114xxU03 ( 855 836 )  100.n
R_D52113LOADxxU03 ( 856 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU03 ( 856 836 )  100.n
R_D52112LOADxxU03 ( 857 0 ) COMPLEX( 3.9963,-2.265)
R_D52112xxU03 ( 857 836 )  100.n
R_D52111LOADxxU03 ( 858 0 ) COMPLEX( 390., 0.)
R_D52111xxU03 ( 858 836 )  1.E+12
R_D52110LOADxxU03 ( 859 0 ) COMPLEX( 8.1777,-4.4139)
R_D52110xxU03 ( 859 836 )  100.n
R_D52109LOADxxU03 ( 860 0 ) COMPLEX( 390., 0.)
R_D52109xxU03 ( 860 836 )  1.E+12
R_D52107xxU03 ( 861 836 )  100.n
R_D52108xxU03 ( 862 836 )  100.n
R_D52108LOADxxU03 ( 0 862 ) COMPLEX( 13.9875,-8.6688)
R_D52107LOADxxU03 ( 0 861 ) COMPLEX( 13.9875,-8.6688)
R_D52106LOADxxU03 ( 0 863 ) COMPLEX( 390., 0.)
R_D52106xxU03 ( 863 836 )  1.E+12
R_D52105LOADxxU03 ( 0 864 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU03 ( 864 836 )  100.n
R_D52104LOADxxU03 ( 0 865 ) COMPLEX( 26.6742,-17.9253)
R_D52104xxU03 ( 865 836 )  100.n
R_D52103LOADxxU03 ( 0 866 ) COMPLEX( 390., 0.)
R_D52103xxU03 ( 866 836 )  1.E+12
R_D52102LOADxxU03 ( 0 867 ) COMPLEX( 390., 0.)
R_D52102xxU03 ( 867 836 )  1.E+12
R_D52101LOADxxU03 ( 0 868 ) COMPLEX( 2.8263,-1.8255)
R_D52101xxU03 ( 836 868 )  100.n
*---------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U04CCM 
R_D52101xxU04 ( 870 902 )  100.n
R_D52101LOADxxU04 ( 0 902 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU04 ( 901 870 )  100.n
R_D52102LOADxxU04 ( 0 901 ) COMPLEX( 390., 0.)
R_D52103xxU04 ( 900 870 )  100.n
R_D52103LOADxxU04 ( 0 900 ) COMPLEX( 390., 0.)
R_D52104xxU04 ( 899 870 )  100.n
R_D52104LOADxxU04 ( 0 899 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU04 ( 898 870 )  100.n
R_D52105LOADxxU04 ( 0 898 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU04 ( 897 870 )  100.n
R_D52106LOADxxU04 ( 0 897 ) COMPLEX( 390., 0.)
R_D52107LOADxxU04 ( 0 895 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU04 ( 0 896 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU04 ( 896 870 )  100.n
R_D52107xxU04 ( 895 870 )  100.n
R_D52109xxU04 ( 894 870 )  100.n
R_D52109LOADxxU04 ( 894 0 ) COMPLEX( 390., 0.)
R_D52110xxU04 ( 893 870 )  100.n
R_D52110LOADxxU04 ( 893 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU04 ( 892 870 )  100.n
R_D52111LOADxxU04 ( 892 0 ) COMPLEX( 390., 0.)
R_D52112xxU04 ( 891 870 )  100.n
R_D52112LOADxxU04 ( 891 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU04 ( 890 870 )  100.n
R_D52113LOADxxU04 ( 890 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU04 ( 889 870 )  100.n
R_D52114LOADxxU04 ( 889 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU04 ( 888 870 )  100.n
R_D52116LOADxxU04 ( 888 0 ) COMPLEX( 390., 0.)
R_D52ExxU04 ( 636 870 )  100.n
R_D52115xxU04 ( 886 870 )  100.n
R_D52115LOADxxU04 ( 886 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU04 ( 870 885 )  100.n
R_D52118LOADxxU04 ( 0 885 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU04 ( 884 870 )  100.n
R_D52119LOADxxU04 ( 0 884 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU04 ( 883 870 )  100.n
R_D52120LOADxxU04 ( 0 883 ) COMPLEX( 390., 0.)
R_D52121xxU04 ( 882 870 )  100.n
R_D52121LOADxxU04 ( 0 882 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU04 ( 881 870 )  100.n
R_D52122LOADxxU04 ( 0 881 ) COMPLEX( 390., 0.)
R_D52123xxU04 ( 880 870 )  100.n
R_D52123LOADxxU04 ( 0 880 ) COMPLEX( 390., 0.)
R_D52124LOADxxU04 ( 0 878 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU04 ( 0 879 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU04 ( 879 870 )  100.n
R_D52124xxU04 ( 878 870 )  100.n
R_D52125xxU04 ( 877 870 )  100.n
R_D52125LOADxxU04 ( 877 0 ) COMPLEX( 390., 0.)
R_D52126xxU04 ( 876 870 )  100.n
R_D52126LOADxxU04 ( 876 0 ) COMPLEX( 390., 0.)
R_D52127xxU04 ( 875 870 )  100.n
R_D52127LOADxxU04 ( 875 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU04 ( 874 870 )  100.n
R_D52128LOADxxU04 ( 874 0 ) COMPLEX( 390., 0.)
R_D52129xxU04 ( 873 870 )  100.n
R_D52129LOADxxU04 ( 873 0 ) COMPLEX( 390., 0.)
R_D52130xxU04 ( 872 870 )  100.n
R_D52130LOADxxU04 ( 872 0 ) COMPLEX( 390., 0.)
R_D52131xxU04 ( 871 870 )  100.n
R_D52131LOADxxU04 ( 871 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU04 ( 869 870 )  100.n
R_D52132LOADxxU04 ( 869 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSSE1 
R_D52E1xxQSSE1 ( 629 905 )  100.n
R_D52E2xxQSSE1 ( 589 909 )  100.n
R_D52307xxQSSE1 ( 918 903 )  100.n
R_D52307LOADxxQSSE1 ( 0 918 ) COMPLEX( 13.9875,-8.6688)
R_D52306xxQSSE1 ( 917 903 )  100.n
R_D52306LOADxxQSSE1 ( 0 917 ) COMPLEX( 390., 0.)
R_D52305xxQSSE1 ( 916 903 )  100.n
R_D52305LOADxxQSSE1 ( 0 916 ) COMPLEX( 390., 0.)
R_D52304xxQSSE1 ( 915 903 )  100.n
R_D52304LOADxxQSSE1 ( 0 915 ) COMPLEX( 13.9875,-8.6688)
R_D52303xxQSSE1 ( 914 903 )  100.n
R_D52303LOADxxQSSE1 ( 0 914 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE1 ( 913 903 )  100.n
R_D52302LOADxxQSSE1 ( 0 913 ) COMPLEX( 26.6742,-17.9253)
R_D52301xxQSSE1 ( 912 903 )  100.n
R_D52301LOADxxQSSE1 ( 0 912 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE1 ( 911 909 )  100.n
R_D52203LOADxxQSSE1 ( 0 911 ) COMPLEX( 390., 0.)
R_D52202xxQSSE1 ( 910 909 )  100.n
R_D52202LOADxxQSSE1 ( 0 910 ) COMPLEX( 390., 0.)
R_D52201xxQSSE1 ( 908 909 )  100.n
R_D52201LOADxxQSSE1 ( 0 908 ) COMPLEX( 17.8179,-11.5092)
R_D52103xxQSSE1 ( 907 905 )  100.n
R_D52103LOADxxQSSE1 ( 0 907 ) COMPLEX( 390., 0.)
R_D52102xxQSSE1 ( 906 905 )  100.n
R_D52102LOADxxQSSE1 ( 0 906 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE1 ( 904 905 )  100.n
R_D52101LOADxxQSSE1 ( 0 904 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE1 ( 0 0 )  1.E+12
R_D52L2xxQSSE1 ( 903 909 )  100.n
*-------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSSE2 
R_D52E1xxQSSE2 ( 581 921 )  100.n
R_D52E2xxQSSE2 ( 638 925 )  100.n
R_D52306xxQSSE2 ( 933 919 )  100.n
R_D52306LOADxxQSSE2 ( 0 933 ) COMPLEX( 390., 0.)
R_D52305xxQSSE2 ( 932 919 )  100.n
R_D52305LOADxxQSSE2 ( 0 932 ) COMPLEX( 390., 0.)
R_D52304xxQSSE2 ( 931 919 )  100.n
R_D52304LOADxxQSSE2 ( 0 931 ) COMPLEX( 390., 0.)
R_D52303xxQSSE2 ( 930 919 )  100.n
R_D52303LOADxxQSSE2 ( 0 930 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE2 ( 929 919 )  100.n
R_D52302LOADxxQSSE2 ( 0 929 ) COMPLEX( 161.6139,-121.2105)
R_D52301xxQSSE2 ( 928 919 )  100.n
R_D52301LOADxxQSSE2 ( 0 928 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE2 ( 927 925 )  100.n
R_D52203LOADxxQSSE2 ( 0 927 ) COMPLEX( 390., 0.)
R_D52202xxQSSE2 ( 926 925 )  100.n
R_D52202LOADxxQSSE2 ( 0 926 ) COMPLEX( 390., 0.)
R_D52201xxQSSE2 ( 924 925 )  100.n
R_D52201LOADxxQSSE2 ( 0 924 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE2 ( 923 921 )  100.n
R_D52103LOADxxQSSE2 ( 0 923 ) COMPLEX( 390., 0.)
R_D52102xxQSSE2 ( 922 921 )  100.n
R_D52102LOADxxQSSE2 ( 0 922 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE2 ( 920 921 )  100.n
R_D52101LOADxxQSSE2 ( 0 920 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE2 ( 0 0 )  1.E+12
R_D52L2xxQSSE2 ( 919 925 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSAM1 
R_D52101xxQSAM1 ( 935 964 )  100.n
R_D52101LOADxxQSAM1 ( 0 964 ) COMPLEX( 26.6742,-17.9253)
R_D52102xxQSAM1 ( 963 935 )  100.n
R_D52102LOADxxQSAM1 ( 0 963 ) COMPLEX( 390., 0.)
R_D52103xxQSAM1 ( 962 935 )  100.n
R_D52103LOADxxQSAM1 ( 0 962 ) COMPLEX( 53.3484,-35.8503)
R_D52104xxQSAM1 ( 961 935 )  100.n
R_D52104LOADxxQSAM1 ( 0 961 ) COMPLEX( 176.6793,-141.7467)
R_D52105xxQSAM1 ( 960 935 )  100.n
R_D52105LOADxxQSAM1 ( 0 960 ) COMPLEX( 390., 0.)
R_D52106xxQSAM1 ( 959 935 )  100.n
R_D52106LOADxxQSAM1 ( 0 959 ) COMPLEX( 26.6742,-17.9253)
R_D52107LOADxxQSAM1 ( 0 958 ) COMPLEX( 23.5224,-11.3925)
R_D52107xxQSAM1 ( 958 935 )  100.n
R_D52108xxQSAM1 ( 957 935 )  100.n
R_D52108LOADxxQSAM1 ( 957 0 ) COMPLEX( 10.4544,-5.0634)
R_D52109xxQSAM1 ( 956 935 )  100.n
R_D52109LOADxxQSAM1 ( 956 0 ) COMPLEX( 390., 0.)
R_D52110xxQSAM1 ( 955 935 )  100.n
R_D52110LOADxxQSAM1 ( 955 0 ) COMPLEX( 71.0055,-49.5621)
R_D52111xxQSAM1 ( 954 935 )  100.n
R_D52111LOADxxQSAM1 ( 954 0 ) COMPLEX( 390., 0.)
R_D52112xxQSAM1 ( 953 935 )  100.n
R_D52112LOADxxQSAM1 ( 953 0 ) COMPLEX( 5.8614,-3.3219)
R_D52113xxQSAM1 ( 952 935 )  100.n
R_D52113LOADxxQSAM1 ( 952 0 ) COMPLEX( 9.7587,-6.048)
R_D52ExxQSAM1 ( 632 935 )  100.n
R_D52114xxQSAM1 ( 950 935 )  100.n
R_D52114LOADxxQSAM1 ( 950 0 ) COMPLEX( 53.3484,-35.8503)
R_D52116xxQSAM1 ( 935 949 )  100.n
R_D52116LOADxxQSAM1 ( 0 949 ) COMPLEX( 9.9912,-6.192)
R_D52117xxQSAM1 ( 948 935 )  100.n
R_D52117LOADxxQSAM1 ( 0 948 ) COMPLEX( 390., 0.)
R_D52118xxQSAM1 ( 947 935 )  100.n
R_D52118LOADxxQSAM1 ( 0 947 ) COMPLEX( 9.9912,-6.192)
R_D52119xxQSAM1 ( 946 935 )  100.n
R_D52119LOADxxQSAM1 ( 0 946 ) COMPLEX( 390., 0.)
R_D52120xxQSAM1 ( 945 935 )  100.n
R_D52120LOADxxQSAM1 ( 0 945 ) COMPLEX( 12.1899,-4.0068)
R_D52121xxQSAM1 ( 944 935 )  100.n
R_D52121LOADxxQSAM1 ( 0 944 ) COMPLEX( 355.0272,-247.8105)
R_D52115LOADxxQSAM1 ( 0 943 ) COMPLEX( 390., 0.)
R_D52115xxQSAM1 ( 943 935 )  100.n
R_D52122xxQSAM1 ( 942 935 )  100.n
R_D52122LOADxxQSAM1 ( 942 0 ) COMPLEX( 13.9875,-8.6688)
R_D52123xxQSAM1 ( 941 935 )  100.n
R_D52123LOADxxQSAM1 ( 941 0 ) COMPLEX( 4.6578,-2.256)
R_D52124xxQSAM1 ( 940 935 )  100.n
R_D52124LOADxxQSAM1 ( 940 0 ) COMPLEX( 39.204,-18.9873)
R_D52125xxQSAM1 ( 939 935 )  100.n
R_D52125LOADxxQSAM1 ( 939 0 ) COMPLEX( 39.204,-18.9873)
R_D52126xxQSAM1 ( 938 935 )  100.n
R_D52126LOADxxQSAM1 ( 938 0 ) COMPLEX( 3.6654,-1.2048)
R_D52127xxQSAM1 ( 937 935 )  100.n
R_D52127LOADxxQSAM1 ( 937 0 ) COMPLEX( 1.1559,-0.5598)
R_D52128xxQSAM1 ( 936 935 )  100.n
R_D52128LOADxxQSAM1 ( 936 0 ) COMPLEX( 1.8093,-0.8763)
R_D52129xxQSAM1 ( 934 935 )  100.n
R_D52129LOADxxQSAM1 ( 934 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSAM2 
R_D52101xxQSAM2 ( 975 991 )  100.n
R_D52101LOADxxQSAM2 ( 0 991 ) COMPLEX( 26.6742,-17.9253)
R_D52102xxQSAM2 ( 990 975 )  100.n
R_D52102LOADxxQSAM2 ( 0 990 ) COMPLEX( 390., 0.)
R_D52103xxQSAM2 ( 989 975 )  100.n
R_D52103LOADxxQSAM2 ( 0 989 ) COMPLEX( 53.3484,-35.8503)
R_D52104xxQSAM2 ( 988 975 )  100.n
R_D52104LOADxxQSAM2 ( 0 988 ) COMPLEX( 176.6793,-141.7467)
R_D52105xxQSAM2 ( 987 975 )  100.n
R_D52105LOADxxQSAM2 ( 0 987 ) COMPLEX( 390., 0.)
R_D52106xxQSAM2 ( 986 975 )  100.n
R_D52106LOADxxQSAM2 ( 0 986 ) COMPLEX( 26.6742,-17.9253)
R_D52107LOADxxQSAM2 ( 0 985 ) COMPLEX( 20.9814,-13.0032)
R_D52107xxQSAM2 ( 985 975 )  100.n
R_D52108xxQSAM2 ( 984 975 )  100.n
R_D52108LOADxxQSAM2 ( 984 0 ) COMPLEX( 9.7692,-5.5365)
R_D52109xxQSAM2 ( 983 975 )  100.n
R_D52109LOADxxQSAM2 ( 983 0 ) COMPLEX( 13.9875,-8.6688)
R_D52110xxQSAM2 ( 982 975 )  100.n
R_D52110LOADxxQSAM2 ( 982 0 ) COMPLEX( 71.0055,-49.5621)
R_D52111xxQSAM2 ( 981 975 )  100.n
R_D52111LOADxxQSAM2 ( 981 0 ) COMPLEX( 390., 0.)
R_D52112xxQSAM2 ( 980 975 )  100.n
R_D52112LOADxxQSAM2 ( 980 0 ) COMPLEX( 5.8614,-3.3219)
R_D52113xxQSAM2 ( 979 975 )  100.n
R_D52113LOADxxQSAM2 ( 979 0 ) COMPLEX( 390., 0.)
R_D52ExxQSAM2 ( 549 975 )  100.n
R_D52114xxQSAM2 ( 977 975 )  100.n
R_D52114LOADxxQSAM2 ( 977 0 ) COMPLEX( 53.3484,-35.8503)
R_D52116xxQSAM2 ( 975 976 )  100.n
R_D52116LOADxxQSAM2 ( 0 976 ) COMPLEX( 390., 0.)
R_D52117xxQSAM2 ( 974 975 )  100.n
R_D52117LOADxxQSAM2 ( 0 974 ) COMPLEX( 390., 0.)
R_D52118xxQSAM2 ( 973 975 )  100.n
R_D52118LOADxxQSAM2 ( 0 973 ) COMPLEX( 390., 0.)
R_D52119xxQSAM2 ( 972 975 )  100.n
R_D52119LOADxxQSAM2 ( 0 972 ) COMPLEX( 390., 0.)
R_D52120xxQSAM2 ( 971 975 )  100.n
R_D52120LOADxxQSAM2 ( 0 971 ) COMPLEX( 390., 0.)
R_D52121xxQSAM2 ( 970 975 )  100.n
R_D52121LOADxxQSAM2 ( 0 970 ) COMPLEX( 235.5726,-188.9955)
R_D52115LOADxxQSAM2 ( 0 969 ) COMPLEX( 390., 0.)
R_D52115xxQSAM2 ( 969 975 )  100.n
R_D52122xxQSAM2 ( 968 975 )  100.n
R_D52122LOADxxQSAM2 ( 968 0 ) COMPLEX( 390., 0.)
R_D52123xxQSAM2 ( 967 975 )  100.n
R_D52123LOADxxQSAM2 ( 967 0 ) COMPLEX( 39.204,-18.9873)
R_D52124xxQSAM2 ( 966 975 )  100.n
R_D52124LOADxxQSAM2 ( 966 0 ) COMPLEX( 39.204,-18.9873)
R_D52125xxQSAM2 ( 965 975 )  100.n
R_D52125LOADxxQSAM2 ( 965 0 ) COMPLEX( 3.6654,-1.2048)
*-------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U05CCM 
R_D52101xxU05 ( 993 1025 )  100.n
R_D52101LOADxxU05 ( 0 1025 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU05 ( 1024 993 )  100.n
R_D52102LOADxxU05 ( 0 1024 ) COMPLEX( 390., 0.)
R_D52103xxU05 ( 1023 993 )  100.n
R_D52103LOADxxU05 ( 0 1023 ) COMPLEX( 390., 0.)
R_D52104xxU05 ( 1022 993 )  100.n
R_D52104LOADxxU05 ( 0 1022 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU05 ( 1021 993 )  100.n
R_D52105LOADxxU05 ( 0 1021 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU05 ( 1020 993 )  100.n
R_D52106LOADxxU05 ( 0 1020 ) COMPLEX( 390., 0.)
R_D52107LOADxxU05 ( 0 1018 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU05 ( 0 1019 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU05 ( 1019 993 )  100.n
R_D52107xxU05 ( 1018 993 )  100.n
R_D52109xxU05 ( 1017 993 )  100.n
R_D52109LOADxxU05 ( 1017 0 ) COMPLEX( 390., 0.)
R_D52110xxU05 ( 1016 993 )  100.n
R_D52110LOADxxU05 ( 1016 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU05 ( 1015 993 )  100.n
R_D52111LOADxxU05 ( 1015 0 ) COMPLEX( 390., 0.)
R_D52112xxU05 ( 1014 993 )  100.n
R_D52112LOADxxU05 ( 1014 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU05 ( 1013 993 )  100.n
R_D52113LOADxxU05 ( 1013 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU05 ( 1012 993 )  100.n
R_D52114LOADxxU05 ( 1012 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU05 ( 1011 993 )  100.n
R_D52116LOADxxU05 ( 1011 0 ) COMPLEX( 390., 0.)
R_D52ExxU05 ( 582 993 )  100.n
R_D52115xxU05 ( 1009 993 )  100.n
R_D52115LOADxxU05 ( 1009 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU05 ( 993 1008 )  100.n
R_D52118LOADxxU05 ( 0 1008 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU05 ( 1007 993 )  100.n
R_D52119LOADxxU05 ( 0 1007 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU05 ( 1006 993 )  100.n
R_D52120LOADxxU05 ( 0 1006 ) COMPLEX( 390., 0.)
R_D52121xxU05 ( 1005 993 )  100.n
R_D52121LOADxxU05 ( 0 1005 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU05 ( 1004 993 )  100.n
R_D52122LOADxxU05 ( 0 1004 ) COMPLEX( 390., 0.)
R_D52123xxU05 ( 1003 993 )  100.n
R_D52123LOADxxU05 ( 0 1003 ) COMPLEX( 390., 0.)
R_D52124LOADxxU05 ( 0 1001 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU05 ( 0 1002 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU05 ( 1002 993 )  100.n
R_D52124xxU05 ( 1001 993 )  100.n
R_D52125xxU05 ( 1000 993 )  100.n
R_D52125LOADxxU05 ( 1000 0 ) COMPLEX( 390., 0.)
R_D52126xxU05 ( 999 993 )  100.n
R_D52126LOADxxU05 ( 999 0 ) COMPLEX( 390., 0.)
R_D52127xxU05 ( 998 993 )  100.n
R_D52127LOADxxU05 ( 998 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU05 ( 997 993 )  100.n
R_D52128LOADxxU05 ( 997 0 ) COMPLEX( 390., 0.)
R_D52129xxU05 ( 996 993 )  100.n
R_D52129LOADxxU05 ( 996 0 ) COMPLEX( 390., 0.)
R_D52130xxU05 ( 995 993 )  100.n
R_D52130LOADxxU05 ( 995 0 ) COMPLEX( 390., 0.)
R_D52131xxU05 ( 994 993 )  100.n
R_D52131LOADxxU05 ( 994 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU05 ( 992 993 )  100.n
R_D52132LOADxxU05 ( 992 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U06CCM 
R_D52101xxU06 ( 1027 1059 )  100.n
R_D52101LOADxxU06 ( 0 1059 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU06 ( 1058 1027 )  100.n
R_D52102LOADxxU06 ( 0 1058 ) COMPLEX( 390., 0.)
R_D52103xxU06 ( 1057 1027 )  100.n
R_D52103LOADxxU06 ( 0 1057 ) COMPLEX( 390., 0.)
R_D52104xxU06 ( 1056 1027 )  100.n
R_D52104LOADxxU06 ( 0 1056 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU06 ( 1055 1027 )  100.n
R_D52105LOADxxU06 ( 0 1055 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU06 ( 1054 1027 )  100.n
R_D52106LOADxxU06 ( 0 1054 ) COMPLEX( 390., 0.)
R_D52107LOADxxU06 ( 0 1052 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU06 ( 0 1053 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU06 ( 1053 1027 )  100.n
R_D52107xxU06 ( 1052 1027 )  100.n
R_D52109xxU06 ( 1051 1027 )  100.n
R_D52109LOADxxU06 ( 1051 0 ) COMPLEX( 390., 0.)
R_D52110xxU06 ( 1050 1027 )  100.n
R_D52110LOADxxU06 ( 1050 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU06 ( 1049 1027 )  100.n
R_D52111LOADxxU06 ( 1049 0 ) COMPLEX( 390., 0.)
R_D52112xxU06 ( 1048 1027 )  100.n
R_D52112LOADxxU06 ( 1048 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU06 ( 1047 1027 )  100.n
R_D52113LOADxxU06 ( 1047 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU06 ( 1046 1027 )  100.n
R_D52114LOADxxU06 ( 1046 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU06 ( 1045 1027 )  100.n
R_D52116LOADxxU06 ( 1045 0 ) COMPLEX( 390., 0.)
R_D52ExxU06 ( 584 1027 )  100.n
R_D52115xxU06 ( 1043 1027 )  100.n
R_D52115LOADxxU06 ( 1043 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU06 ( 1027 1042 )  100.n
R_D52118LOADxxU06 ( 0 1042 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU06 ( 1041 1027 )  100.n
R_D52119LOADxxU06 ( 0 1041 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU06 ( 1040 1027 )  100.n
R_D52120LOADxxU06 ( 0 1040 ) COMPLEX( 390., 0.)
R_D52121xxU06 ( 1039 1027 )  100.n
R_D52121LOADxxU06 ( 0 1039 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU06 ( 1038 1027 )  100.n
R_D52122LOADxxU06 ( 0 1038 ) COMPLEX( 390., 0.)
R_D52123xxU06 ( 1037 1027 )  100.n
R_D52123LOADxxU06 ( 0 1037 ) COMPLEX( 390., 0.)
R_D52124LOADxxU06 ( 0 1035 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU06 ( 0 1036 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU06 ( 1036 1027 )  100.n
R_D52124xxU06 ( 1035 1027 )  100.n
R_D52125xxU06 ( 1034 1027 )  100.n
R_D52125LOADxxU06 ( 1034 0 ) COMPLEX( 390., 0.)
R_D52126xxU06 ( 1033 1027 )  100.n
R_D52126LOADxxU06 ( 1033 0 ) COMPLEX( 390., 0.)
R_D52127xxU06 ( 1032 1027 )  100.n
R_D52127LOADxxU06 ( 1032 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU06 ( 1031 1027 )  100.n
R_D52128LOADxxU06 ( 1031 0 ) COMPLEX( 390., 0.)
R_D52129xxU06 ( 1030 1027 )  100.n
R_D52129LOADxxU06 ( 1030 0 ) COMPLEX( 390., 0.)
R_D52130xxU06 ( 1029 1027 )  100.n
R_D52130LOADxxU06 ( 1029 0 ) COMPLEX( 390., 0.)
R_D52131xxU06 ( 1028 1027 )  100.n
R_D52131LOADxxU06 ( 1028 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU06 ( 1026 1027 )  100.n
R_D52132LOADxxU06 ( 1026 0 ) COMPLEX( 390., 0.)
*-------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U07CCM 
R_D52101xxU07 ( 1061 1093 )  100.n
R_D52101LOADxxU07 ( 0 1093 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU07 ( 1092 1061 )  100.n
R_D52102LOADxxU07 ( 0 1092 ) COMPLEX( 390., 0.)
R_D52103xxU07 ( 1091 1061 )  100.n
R_D52103LOADxxU07 ( 0 1091 ) COMPLEX( 390., 0.)
R_D52104xxU07 ( 1090 1061 )  100.n
R_D52104LOADxxU07 ( 0 1090 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU07 ( 1089 1061 )  100.n
R_D52105LOADxxU07 ( 0 1089 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU07 ( 1088 1061 )  100.n
R_D52106LOADxxU07 ( 0 1088 ) COMPLEX( 390., 0.)
R_D52107LOADxxU07 ( 0 1086 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU07 ( 0 1087 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU07 ( 1087 1061 )  100.n
R_D52107xxU07 ( 1086 1061 )  100.n
R_D52109xxU07 ( 1085 1061 )  100.n
R_D52109LOADxxU07 ( 1085 0 ) COMPLEX( 390., 0.)
R_D52110xxU07 ( 1084 1061 )  100.n
R_D52110LOADxxU07 ( 1084 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU07 ( 1083 1061 )  100.n
R_D52111LOADxxU07 ( 1083 0 ) COMPLEX( 390., 0.)
R_D52112xxU07 ( 1082 1061 )  100.n
R_D52112LOADxxU07 ( 1082 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU07 ( 1081 1061 )  100.n
R_D52113LOADxxU07 ( 1081 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU07 ( 1080 1061 )  100.n
R_D52114LOADxxU07 ( 1080 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU07 ( 1079 1061 )  100.n
R_D52116LOADxxU07 ( 1079 0 ) COMPLEX( 390., 0.)
R_D52ExxU07 ( 588 1061 )  100.n
R_D52115xxU07 ( 1077 1061 )  100.n
R_D52115LOADxxU07 ( 1077 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU07 ( 1061 1076 )  100.n
R_D52118LOADxxU07 ( 0 1076 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU07 ( 1075 1061 )  100.n
R_D52119LOADxxU07 ( 0 1075 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU07 ( 1074 1061 )  100.n
R_D52120LOADxxU07 ( 0 1074 ) COMPLEX( 390., 0.)
R_D52121xxU07 ( 1073 1061 )  100.n
R_D52121LOADxxU07 ( 0 1073 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU07 ( 1072 1061 )  100.n
R_D52122LOADxxU07 ( 0 1072 ) COMPLEX( 390., 0.)
R_D52123xxU07 ( 1071 1061 )  100.n
R_D52123LOADxxU07 ( 0 1071 ) COMPLEX( 390., 0.)
R_D52124LOADxxU07 ( 0 1069 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU07 ( 0 1070 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU07 ( 1070 1061 )  100.n
R_D52124xxU07 ( 1069 1061 )  100.n
R_D52125xxU07 ( 1068 1061 )  100.n
R_D52125LOADxxU07 ( 1068 0 ) COMPLEX( 390., 0.)
R_D52126xxU07 ( 1067 1061 )  100.n
R_D52126LOADxxU07 ( 1067 0 ) COMPLEX( 390., 0.)
R_D52127xxU07 ( 1066 1061 )  100.n
R_D52127LOADxxU07 ( 1066 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU07 ( 1065 1061 )  100.n
R_D52128LOADxxU07 ( 1065 0 ) COMPLEX( 390., 0.)
R_D52129xxU07 ( 1064 1061 )  100.n
R_D52129LOADxxU07 ( 1064 0 ) COMPLEX( 390., 0.)
R_D52130xxU07 ( 1063 1061 )  100.n
R_D52130LOADxxU07 ( 1063 0 ) COMPLEX( 390., 0.)
R_D52131xxU07 ( 1062 1061 )  100.n
R_D52131LOADxxU07 ( 1062 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU07 ( 1060 1061 )  100.n
R_D52132LOADxxU07 ( 1060 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U08CCM 
R_D52101xxU08 ( 1095 1127 )  100.n
R_D52101LOADxxU08 ( 0 1127 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU08 ( 1126 1095 )  100.n
R_D52102LOADxxU08 ( 0 1126 ) COMPLEX( 390., 0.)
R_D52103xxU08 ( 1125 1095 )  100.n
R_D52103LOADxxU08 ( 0 1125 ) COMPLEX( 390., 0.)
R_D52104xxU08 ( 1124 1095 )  100.n
R_D52104LOADxxU08 ( 0 1124 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU08 ( 1123 1095 )  100.n
R_D52105LOADxxU08 ( 0 1123 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU08 ( 1122 1095 )  100.n
R_D52106LOADxxU08 ( 0 1122 ) COMPLEX( 390., 0.)
R_D52107LOADxxU08 ( 0 1120 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU08 ( 0 1121 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU08 ( 1121 1095 )  100.n
R_D52107xxU08 ( 1120 1095 )  100.n
R_D52109xxU08 ( 1119 1095 )  100.n
R_D52109LOADxxU08 ( 1119 0 ) COMPLEX( 390., 0.)
R_D52110xxU08 ( 1118 1095 )  100.n
R_D52110LOADxxU08 ( 1118 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU08 ( 1117 1095 )  100.n
R_D52111LOADxxU08 ( 1117 0 ) COMPLEX( 390., 0.)
R_D52112xxU08 ( 1116 1095 )  100.n
R_D52112LOADxxU08 ( 1116 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU08 ( 1115 1095 )  100.n
R_D52113LOADxxU08 ( 1115 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU08 ( 1114 1095 )  100.n
R_D52114LOADxxU08 ( 1114 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU08 ( 1113 1095 )  100.n
R_D52116LOADxxU08 ( 1113 0 ) COMPLEX( 390., 0.)
R_D52ExxU08 ( 587 1095 )  100.n
R_D52115xxU08 ( 1111 1095 )  100.n
R_D52115LOADxxU08 ( 1111 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU08 ( 1095 1110 )  100.n
R_D52118LOADxxU08 ( 0 1110 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU08 ( 1109 1095 )  100.n
R_D52119LOADxxU08 ( 0 1109 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU08 ( 1108 1095 )  100.n
R_D52120LOADxxU08 ( 0 1108 ) COMPLEX( 390., 0.)
R_D52121xxU08 ( 1107 1095 )  100.n
R_D52121LOADxxU08 ( 0 1107 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU08 ( 1106 1095 )  100.n
R_D52122LOADxxU08 ( 0 1106 ) COMPLEX( 390., 0.)
R_D52123xxU08 ( 1105 1095 )  100.n
R_D52123LOADxxU08 ( 0 1105 ) COMPLEX( 390., 0.)
R_D52124LOADxxU08 ( 0 1103 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU08 ( 0 1104 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU08 ( 1104 1095 )  100.n
R_D52124xxU08 ( 1103 1095 )  100.n
R_D52125xxU08 ( 1102 1095 )  100.n
R_D52125LOADxxU08 ( 1102 0 ) COMPLEX( 390., 0.)
R_D52126xxU08 ( 1101 1095 )  100.n
R_D52126LOADxxU08 ( 1101 0 ) COMPLEX( 390., 0.)
R_D52127xxU08 ( 1100 1095 )  100.n
R_D52127LOADxxU08 ( 1100 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU08 ( 1099 1095 )  100.n
R_D52128LOADxxU08 ( 1099 0 ) COMPLEX( 390., 0.)
R_D52129xxU08 ( 1098 1095 )  100.n
R_D52129LOADxxU08 ( 1098 0 ) COMPLEX( 390., 0.)
R_D52130xxU08 ( 1097 1095 )  100.n
R_D52130LOADxxU08 ( 1097 0 ) COMPLEX( 390., 0.)
R_D52131xxU08 ( 1096 1095 )  100.n
R_D52131LOADxxU08 ( 1096 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU08 ( 1094 1095 )  100.n
R_D52132LOADxxU08 ( 1094 0 ) COMPLEX( 390., 0.)
*---------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA CCME1 
R_D52E1xxCCME1 ( 583 1129 )  100.n
R_D52E2xxCCME1 ( 597 1128 )  100.n
R_D52206xxCCME1 ( 1142 1128 )  100.n
R_D52206LOADxxCCME1 ( 0 1142 ) COMPLEX( 390., 0.)
R_D52205xxCCME1 ( 1141 1128 )  100.n
R_D52205LOADxxCCME1 ( 0 1141 ) COMPLEX( 390., 0.)
R_D52204xxCCME1 ( 1140 1128 )  100.n
R_D52204LOADxxCCME1 ( 0 1140 ) COMPLEX( 390., 0.)
R_D52203xxCCME1 ( 1139 1128 )  100.n
R_D52203LOADxxCCME1 ( 0 1139 ) COMPLEX( 390., 0.)
R_D52202xxCCME1 ( 1138 1128 )  100.n
R_D52202LOADxxCCME1 ( 0 1138 ) COMPLEX( 3.9963,-2.265)
R_D52201xxCCME1 ( 1137 1128 )  100.n
R_D52201LOADxxCCME1 ( 0 1137 ) COMPLEX( 3.9963,-2.265)
R_D52107xxCCME1 ( 1136 1129 )  100.n
R_D52107LOADxxCCME1 ( 0 1136 ) COMPLEX( 1.363267K,-1.593835K)
R_D52106xxCCME1 ( 1135 1129 )  100.n
R_D52106LOADxxCCME1 ( 0 1135 ) COMPLEX( 390., 0.)
R_D52105xxCCME1 ( 1134 1129 )  100.n
R_D52105LOADxxCCME1 ( 0 1134 ) COMPLEX( 30.976, 0.)
R_D52104xxCCME1 ( 1133 1129 )  100.n
R_D52104LOADxxCCME1 ( 0 1133 ) COMPLEX( 33.3429,-22.4064)
R_D52103xxCCME1 ( 1132 1129 )  100.n
R_D52103LOADxxCCME1 ( 0 1132 ) COMPLEX( 390., 0.)
R_D52102xxCCME1 ( 1131 1129 )  100.n
R_D52102LOADxxCCME1 ( 0 1131 ) COMPLEX( 3.9963,-2.265)
R_D52101xxCCME1 ( 1130 1129 )  100.n
R_D52101LOADxxCCME1 ( 0 1130 ) COMPLEX( 2.97,-2.6193)
R_D52LxxCCME1 ( 0 0 )  1.E+12
*------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA CCME2 
R_D52E1xxCCME2 ( 572 1144 )  100.n
R_D52E2xxCCME2 ( 565 1143 )  100.n
R_D52206xxCCME2 ( 1157 1143 )  100.n
R_D52206LOADxxCCME2 ( 0 1157 ) COMPLEX( 390., 0.)
R_D52205xxCCME2 ( 1156 1143 )  100.n
R_D52205LOADxxCCME2 ( 0 1156 ) COMPLEX( 390., 0.)
R_D52204xxCCME2 ( 1155 1143 )  100.n
R_D52204LOADxxCCME2 ( 0 1155 ) COMPLEX( 390., 0.)
R_D52203xxCCME2 ( 1154 1143 )  100.n
R_D52203LOADxxCCME2 ( 0 1154 ) COMPLEX( 390., 0.)
R_D52202xxCCME2 ( 1153 1143 )  100.n
R_D52202LOADxxCCME2 ( 0 1153 ) COMPLEX( 3.9963,-2.265)
R_D52201xxCCME2 ( 1152 1143 )  100.n
R_D52201LOADxxCCME2 ( 0 1152 ) COMPLEX( 3.9963,-2.265)
R_D52107xxCCME2 ( 1151 1144 )  100.n
R_D52107LOADxxCCME2 ( 0 1151 ) COMPLEX( 1.363267K,-1.593835K)
R_D52106xxCCME2 ( 1150 1144 )  100.n
R_D52106LOADxxCCME2 ( 0 1150 ) COMPLEX( 390., 0.)
R_D52105xxCCME2 ( 1149 1144 )  100.n
R_D52105LOADxxCCME2 ( 0 1149 ) COMPLEX( 30.976, 0.)
R_D52104xxCCME2 ( 1148 1144 )  100.n
R_D52104LOADxxCCME2 ( 0 1148 ) COMPLEX( 33.3429,-22.4064)
R_D52103xxCCME2 ( 1147 1144 )  100.n
R_D52103LOADxxCCME2 ( 0 1147 ) COMPLEX( 390., 0.)
R_D52102xxCCME2 ( 1146 1144 )  100.n
R_D52102LOADxxCCME2 ( 0 1146 ) COMPLEX( 3.9963,-2.265)
R_D52101xxCCME2 ( 1145 1144 )  100.n
R_D52101LOADxxCCME2 ( 0 1145 ) COMPLEX( 2.97,-2.6193)
R_D52LxxCCME2 ( 0 0 )  1.E+12
*---------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA CCMD1 
R_D52101xxCCMD1 ( 1180 1159 )  100.n
R_D52101LOADxxCCMD1 ( 0 1180 ) COMPLEX( 168.96,-126.72)
R_D52E1xxCCMD1 ( 454 1159 )  100.n
R_D52209xxCCMD1 ( 1178 1169 )  100.n
R_D52209LOADxxCCMD1 ( 0 1178 ) COMPLEX( 390., 0.)
R_D52E2xxCCMD1 ( 595 1169 )  100.n
R_D52208xxCCMD1 ( 1176 1169 )  100.n
R_D52208LOADxxCCMD1 ( 0 1176 ) COMPLEX( 1.363267K,-1.593835K)
R_D52207xxCCMD1 ( 1175 1169 )  100.n
R_D52207LOADxxCCMD1 ( 0 1175 ) COMPLEX( 235.5726,-188.9955)
R_D52206xxCCMD1 ( 1174 1169 )  100.n
R_D52206LOADxxCCMD1 ( 0 1174 ) COMPLEX( 5.8614,-3.3219)
R_D52205xxCCMD1 ( 1173 1169 )  100.n
R_D52205LOADxxCCMD1 ( 0 1173 ) COMPLEX( 11.6097,-6.8889)
R_D52204xxCCMD1 ( 1172 1169 )  100.n
R_D52204LOADxxCCMD1 ( 0 1172 ) COMPLEX( 390., 0.)
R_D52203xxCCMD1 ( 1171 1169 )  100.n
R_D52203LOADxxCCMD1 ( 0 1171 ) COMPLEX( 1.363267K,-1.593835K)
R_D52202xxCCMD1 ( 1170 1169 )  100.n
R_D52202LOADxxCCMD1 ( 0 1170 ) COMPLEX( 235.5726,-188.9955)
R_D52201xxCCMD1 ( 1168 1169 )  100.n
R_D52201LOADxxCCMD1 ( 0 1168 ) COMPLEX( 168.96,-126.72)
R_D52110xxCCMD1 ( 1167 1159 )  100.n
R_D52110LOADxxCCMD1 ( 0 1167 ) COMPLEX( 390., 0.)
R_D52109xxCCMD1 ( 1166 1159 )  100.n
R_D52109LOADxxCCMD1 ( 0 1166 ) COMPLEX( 11.6097,-6.8889)
R_D52108xxCCMD1 ( 1165 1159 )  100.n
R_D52108LOADxxCCMD1 ( 0 1165 ) COMPLEX( 11.6097,-6.8889)
R_D52107xxCCMD1 ( 1164 1159 )  100.n
R_D52107LOADxxCCMD1 ( 0 1164 ) COMPLEX( 390., 0.)
R_D52106xxCCMD1 ( 1163 1159 )  100.n
R_D52106LOADxxCCMD1 ( 0 1163 ) COMPLEX( 390., 0.)
R_D52105xxCCMD1 ( 1162 1159 )  100.n
R_D52105LOADxxCCMD1 ( 0 1162 ) COMPLEX( 5.8614,-3.3219)
R_D52104xxCCMD1 ( 1161 1159 )  100.n
R_D52104LOADxxCCMD1 ( 0 1161 ) COMPLEX( 5.8614,-3.3219)
R_D52103xxCCMD1 ( 1160 1159 )  100.n
R_D52103LOADxxCCMD1 ( 0 1160 ) COMPLEX( 390., 0.)
R_D52102xxCCMD1 ( 1158 1159 )  100.n
R_D52102LOADxxCCMD1 ( 0 1158 ) COMPLEX( 1.363267K,-1.593835K)
R_D52LxxCCMD1 ( 0 0 )  1.E+12
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA CCMD2 
R_D52101xxCCMD2 ( 1203 1182 )  100.n
R_D52101LOADxxCCMD2 ( 0 1203 ) COMPLEX( 168.96,-126.72)
R_D52E1xxCCMD2 ( 567 1182 )  100.n
R_D52209xxCCMD2 ( 1201 1192 )  100.n
R_D52209LOADxxCCMD2 ( 0 1201 ) COMPLEX( 390., 0.)
R_D52E2xxCCMD2 ( 560 1192 )  100.n
R_D52208xxCCMD2 ( 1199 1192 )  100.n
R_D52208LOADxxCCMD2 ( 0 1199 ) COMPLEX( 1.363267K,-1.593835K)
R_D52207xxCCMD2 ( 1198 1192 )  100.n
R_D52207LOADxxCCMD2 ( 0 1198 ) COMPLEX( 235.5726,-188.9955)
R_D52206xxCCMD2 ( 1197 1192 )  100.n
R_D52206LOADxxCCMD2 ( 0 1197 ) COMPLEX( 5.8614,-3.3219)
R_D52205xxCCMD2 ( 1196 1192 )  100.n
R_D52205LOADxxCCMD2 ( 0 1196 ) COMPLEX( 11.6097,-6.8889)
R_D52204xxCCMD2 ( 1195 1192 )  100.n
R_D52204LOADxxCCMD2 ( 0 1195 ) COMPLEX( 390., 0.)
R_D52203xxCCMD2 ( 1194 1192 )  100.n
R_D52203LOADxxCCMD2 ( 0 1194 ) COMPLEX( 1.363267K,-1.593835K)
R_D52202xxCCMD2 ( 1193 1192 )  100.n
R_D52202LOADxxCCMD2 ( 0 1193 ) COMPLEX( 235.5726,-188.9955)
R_D52201xxCCMD2 ( 1191 1192 )  100.n
R_D52201LOADxxCCMD2 ( 0 1191 ) COMPLEX( 168.96,-126.72)
R_D52110xxCCMD2 ( 1190 1182 )  100.n
R_D52110LOADxxCCMD2 ( 0 1190 ) COMPLEX( 390., 0.)
R_D52109xxCCMD2 ( 1189 1182 )  100.n
R_D52109LOADxxCCMD2 ( 0 1189 ) COMPLEX( 11.6097,-6.8889)
R_D52108xxCCMD2 ( 1188 1182 )  100.n
R_D52108LOADxxCCMD2 ( 0 1188 ) COMPLEX( 11.6097,-6.8889)
R_D52107xxCCMD2 ( 1187 1182 )  100.n
R_D52107LOADxxCCMD2 ( 0 1187 ) COMPLEX( 390., 0.)
R_D52106xxCCMD2 ( 1186 1182 )  100.n
R_D52106LOADxxCCMD2 ( 0 1186 ) COMPLEX( 390., 0.)
R_D52105xxCCMD2 ( 1185 1182 )  100.n
R_D52105LOADxxCCMD2 ( 0 1185 ) COMPLEX( 5.8614,-3.3219)
R_D52104xxCCMD2 ( 1184 1182 )  100.n
R_D52104LOADxxCCMD2 ( 0 1184 ) COMPLEX( 5.8614,-3.3219)
R_D52103xxCCMD2 ( 1183 1182 )  100.n
R_D52103LOADxxCCMD2 ( 0 1183 ) COMPLEX( 390., 0.)
R_D52102xxCCMD2 ( 1181 1182 )  100.n
R_D52102LOADxxCCMD2 ( 0 1181 ) COMPLEX( 1.363267K,-1.593835K)
R_D52LxxCCMD2 ( 0 0 )  1.E+12
*----------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSSE3 
R_D52E1xxQSSE3 ( 593 1206 )  100.n
R_D52E2xxQSSE3 ( 622 1209 )  100.n
R_D52307xxQSSE3 ( 1218 1204 )  100.n
R_D52307LOADxxQSSE3 ( 0 1218 ) COMPLEX( 390., 0.)
R_D52306xxQSSE3 ( 1217 1204 )  100.n
R_D52306LOADxxQSSE3 ( 0 1217 ) COMPLEX( 390., 0.)
R_D52305xxQSSE3 ( 1216 1204 )  100.n
R_D52305LOADxxQSSE3 ( 0 1216 ) COMPLEX( 390., 0.)
R_D52304xxQSSE3 ( 1215 1204 )  100.n
R_D52304LOADxxQSSE3 ( 0 1215 ) COMPLEX( 390., 0.)
R_D52303xxQSSE3 ( 1214 1204 )  100.n
R_D52303LOADxxQSSE3 ( 0 1214 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE3 ( 1213 1204 )  100.n
R_D52302LOADxxQSSE3 ( 0 1213 ) COMPLEX( 26.6742,-17.9253)
R_D52301xxQSSE3 ( 1212 1204 )  100.n
R_D52301LOADxxQSSE3 ( 0 1212 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE3 ( 1211 1209 )  100.n
R_D52203LOADxxQSSE3 ( 0 1211 ) COMPLEX( 390., 0.)
R_D52202xxQSSE3 ( 1210 1209 )  100.n
R_D52202LOADxxQSSE3 ( 0 1210 ) COMPLEX( 390., 0.)
R_D52201xxQSSE3 ( 1208 1209 )  100.n
R_D52201LOADxxQSSE3 ( 0 1208 ) COMPLEX( 30.976, 0.)
R_D52102xxQSSE3 ( 1207 1206 )  100.n
R_D52102LOADxxQSSE3 ( 0 1207 ) COMPLEX( 30.976, 0.)
R_D52101xxQSSE3 ( 1205 1206 )  100.n
R_D52101LOADxxQSSE3 ( 0 1205 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE3 ( 0 0 )  1.E+12
R_D52L2xxQSSE3 ( 1204 1209 )  100.n
*------------------------------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA QSSE4 
R_D52E1xxQSSE4 ( 616 1221 )  100.n
R_D52E2xxQSSE4 ( 601 1225 )  100.n
R_D52307xxQSSE4 ( 1234 1219 )  100.n
R_D52307LOADxxQSSE4 ( 0 1234 ) COMPLEX( 390., 0.)
R_D52306xxQSSE4 ( 1233 1219 )  100.n
R_D52306LOADxxQSSE4 ( 0 1233 ) COMPLEX( 390., 0.)
R_D52305xxQSSE4 ( 1232 1219 )  100.n
R_D52305LOADxxQSSE4 ( 0 1232 ) COMPLEX( 390., 0.)
R_D52304xxQSSE4 ( 1231 1219 )  100.n
R_D52304LOADxxQSSE4 ( 0 1231 ) COMPLEX( 13.9875,-8.6688)
R_D52303xxQSSE4 ( 1230 1219 )  100.n
R_D52303LOADxxQSSE4 ( 0 1230 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE4 ( 1229 1219 )  100.n
R_D52302LOADxxQSSE4 ( 0 1229 ) COMPLEX( 26.6742,-17.9253)
R_D52301xxQSSE4 ( 1228 1219 )  100.n
R_D52301LOADxxQSSE4 ( 0 1228 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE4 ( 1227 1225 )  100.n
R_D52203LOADxxQSSE4 ( 0 1227 ) COMPLEX( 390., 0.)
R_D52202xxQSSE4 ( 1226 1225 )  100.n
R_D52202LOADxxQSSE4 ( 0 1226 ) COMPLEX( 390., 0.)
R_D52201xxQSSE4 ( 1224 1225 )  100.n
R_D52201LOADxxQSSE4 ( 0 1224 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE4 ( 1223 1221 )  100.n
R_D52103LOADxxQSSE4 ( 0 1223 ) COMPLEX( 390., 0.)
R_D52102xxQSSE4 ( 1222 1221 )  100.n
R_D52102LOADxxQSSE4 ( 0 1222 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE4 ( 1220 1221 )  100.n
R_D52101LOADxxQSSE4 ( 0 1220 ) COMPLEX( 390., 0.)
R_D52L1xxQSSE4 ( 0 0 )  1.E+12
R_D52L2xxQSSE4 ( 1219 1225 )  100.n
*-------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSG3 
R_D52101xxQSG3 ( 1241 1301 )  100.n
R_D52101LOADxxQSG3 ( 0 1301 ) COMPLEX( 390., 0.)
R_D52102xxQSG3 ( 1300 1241 )  100.n
R_D52102LOADxxQSG3 ( 0 1300 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG3 ( 1299 1241 )  100.n
R_D52103LOADxxQSG3 ( 0 1299 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG3 ( 1298 1241 )  100.n
R_D52104LOADxxQSG3 ( 0 1298 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG3 ( 1297 1241 )  100.n
R_D52105LOADxxQSG3 ( 0 1297 ) COMPLEX( 390., 0.)
R_D52107xxQSG3 ( 1296 1241 )  100.n
R_D52107LOADxxQSG3 ( 0 1296 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG3 ( 0 1295 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG3 ( 1295 1241 )  100.n
R_D52110xxQSG3 ( 1294 1241 )  100.n
R_D52110LOADxxQSG3 ( 1294 0 ) COMPLEX( 390., 0.)
R_D52111xxQSG3 ( 1293 1241 )  100.n
R_D52111LOADxxQSG3 ( 1293 0 ) COMPLEX( 16.3926,-10.5885)
R_D52112xxQSG3 ( 1292 1241 )  100.n
R_D52112LOADxxQSG3 ( 1292 0 ) COMPLEX( 235.5726,-188.9955)
R_D52113xxQSG3 ( 1291 1241 )  100.n
R_D52113LOADxxQSG3 ( 1291 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG3 ( 1290 1241 )  100.n
R_D52114LOADxxQSG3 ( 1290 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG3 ( 1289 1241 )  100.n
R_D52115LOADxxQSG3 ( 1289 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG3 ( 0 0 )  1.E+12
R_D52116xxQSG3 ( 1287 1241 )  100.n
R_D52116LOADxxQSG3 ( 1287 0 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG3 ( 1286 1241 )  100.n
R_D52109LOADxxQSG3 ( 1286 0 ) COMPLEX( 3.9963,-2.265)
R_D52L2xxQSG3 ( 1236 1267 )  100.n
R_D52E2xxQSG3 ( 618 1267 )  100.n
R_D52E1xxQSG3 ( 592 1241 )  100.n
R_D52201xxQSG3 ( 1267 1284 )  100.n
R_D52201LOADxxQSG3 ( 0 1284 ) COMPLEX( 390., 0.)
R_D52202xxQSG3 ( 1283 1267 )  100.n
R_D52202LOADxxQSG3 ( 0 1283 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG3 ( 1282 1267 )  100.n
R_D52203LOADxxQSG3 ( 0 1282 ) COMPLEX( 30.976, 0.)
R_D52204xxQSG3 ( 1281 1267 )  100.n
R_D52204LOADxxQSG3 ( 0 1281 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG3 ( 1280 1267 )  100.n
R_D52205LOADxxQSG3 ( 0 1280 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG3 ( 1279 1267 )  100.n
R_D52206LOADxxQSG3 ( 0 0 )  1.E+12
R_D52208LOADxxQSG3 ( 0 1278 ) COMPLEX( 390., 0.)
R_D52208xxQSG3 ( 1278 1267 )  100.n
R_D52210xxQSG3 ( 1277 1267 )  100.n
R_D52210LOADxxQSG3 ( 1277 0 ) COMPLEX( 390., 0.)
R_D52211xxQSG3 ( 1276 1267 )  100.n
R_D52211LOADxxQSG3 ( 1276 0 ) COMPLEX( 123.9039,-92.928)
R_D52212xxQSG3 ( 1275 1267 )  100.n
R_D52212LOADxxQSG3 ( 1275 0 ) COMPLEX( 390., 0.)
R_D52213xxQSG3 ( 1274 1267 )  100.n
R_D52213LOADxxQSG3 ( 1274 0 ) COMPLEX( 235.5726,-188.9955)
R_D52214xxQSG3 ( 1273 1267 )  100.n
R_D52214LOADxxQSG3 ( 1273 0 ) COMPLEX( 168.96,-126.72)
R_D52215xxQSG3 ( 1272 1267 )  100.n
R_D52215LOADxxQSG3 ( 1272 0 ) COMPLEX( 390., 0.)
R_D52216xxQSG3 ( 1271 1267 )  100.n
R_D52216LOADxxQSG3 ( 1271 0 ) COMPLEX( 3.9963,-2.265)
R_D52209xxQSG3 ( 1270 1267 )  100.n
R_D52209LOADxxQSG3 ( 1270 0 ) COMPLEX( 390., 0.)
R_D52326xxQSG3 ( 1269 1236 )  100.n
R_D52326LOADxxQSG3 ( 1269 0 ) COMPLEX( 6.078,-3.2805)
R_D52327xxQSG3 ( 1268 1236 )  100.n
R_D52327LOADxxQSG3 ( 1268 0 ) COMPLEX( 20.4906,-13.2357)
R_D52207LOADxxQSG3 ( 1266 0 ) COMPLEX( 390., 0.)
R_D52207xxQSG3 ( 1266 1267 )  100.n
R_D52301xxQSG3 ( 1236 1264 )  100.n
R_D52301LOADxxQSG3 ( 0 1264 ) COMPLEX( 2.0445,-1.1034)
R_D52302xxQSG3 ( 1263 1236 )  100.n
R_D52302LOADxxQSG3 ( 0 1263 ) COMPLEX( 390., 0.)
R_D52303xxQSG3 ( 1262 1236 )  100.n
R_D52303LOADxxQSG3 ( 0 1262 ) COMPLEX( 176.6793,-141.7467)
R_D52304xxQSG3 ( 1261 1236 )  100.n
R_D52304LOADxxQSG3 ( 0 1261 ) COMPLEX( 390., 0.)
R_D52305xxQSG3 ( 1260 1236 )  100.n
R_D52305LOADxxQSG3 ( 0 1260 ) COMPLEX( 390., 0.)
R_D52306xxQSG3 ( 1259 1236 )  100.n
R_D52306LOADxxQSG3 ( 0 1259 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG3 ( 0 1258 ) COMPLEX( 64.2471,-51.5442)
R_D52308xxQSG3 ( 1258 1236 )  100.n
R_D52311xxQSG3 ( 1257 1236 )  100.n
R_D52311LOADxxQSG3 ( 1257 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG3 ( 1256 1236 )  100.n
R_D52312LOADxxQSG3 ( 1256 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG3 ( 1255 1236 )  100.n
R_D52313LOADxxQSG3 ( 1255 0 ) COMPLEX( 168.96,-126.72)
R_D52314xxQSG3 ( 1254 1236 )  100.n
R_D52314LOADxxQSG3 ( 1254 0 ) COMPLEX( 355.0272,-247.8105)
R_D52315xxQSG3 ( 1253 1236 )  100.n
R_D52315LOADxxQSG3 ( 1253 0 ) COMPLEX( 390., 0.)
R_D52316xxQSG3 ( 1252 1236 )  100.n
R_D52316LOADxxQSG3 ( 1252 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG3 ( 1251 1236 )  100.n
R_D52317LOADxxQSG3 ( 1251 0 ) COMPLEX( 390., 0.)
R_D52310xxQSG3 ( 1250 1236 )  100.n
R_D52310LOADxxQSG3 ( 1250 0 ) COMPLEX( 390., 0.)
R_D52318xxQSG3 ( 1249 1236 )  100.n
R_D52318LOADxxQSG3 ( 1249 0 ) COMPLEX( 390., 0.)
R_D52319xxQSG3 ( 1248 1236 )  100.n
R_D52319LOADxxQSG3 ( 1248 0 ) COMPLEX( 390., 0.)
R_D52309LOADxxQSG3 ( 0 1247 ) COMPLEX( 390., 0.)
R_D52309xxQSG3 ( 1247 1236 )  100.n
R_D52307LOADxxQSG3 ( 1246 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG3 ( 1246 1236 )  100.n
R_D52320xxQSG3 ( 1236 1245 )  100.n
R_D52320LOADxxQSG3 ( 0 1245 ) COMPLEX( 20.4906,-13.2357)
R_D52321xxQSG3 ( 1244 1236 )  100.n
R_D52321LOADxxQSG3 ( 0 1244 ) COMPLEX( 5.8614,-3.3219)
R_D52325xxQSG3 ( 1243 1236 )  100.n
R_D52325LOADxxQSG3 ( 1243 0 ) COMPLEX( 6.078,-3.2805)
R_D52324xxQSG3 ( 1242 1236 )  100.n
R_D52324LOADxxQSG3 ( 1242 0 ) COMPLEX( 32.1234,-25.7721)
R_D52106LOADxxQSG3 ( 0 0 )  1.E+12
R_D52106xxQSG3 ( 1240 1241 )  100.n
R_D52322xxQSG3 ( 1238 1236 )  100.n
R_D52322LOADxxQSG3 ( 0 1238 ) COMPLEX( 5.8614,-3.3219)
R_D52323xxQSG3 ( 1237 1236 )  100.n
R_D52323LOADxxQSG3 ( 0 1237 ) COMPLEX( 390., 0.)
R_D52328xxQSG3 ( 1235 1236 )  100.n
R_D52328LOADxxQSG3 ( 1235 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG4 
R_D52101xxQSG4 ( 1346 1361 )  100.n
R_D52101LOADxxQSG4 ( 0 1361 ) COMPLEX( 390., 0.)
R_D52102xxQSG4 ( 1360 1346 )  100.n
R_D52102LOADxxQSG4 ( 0 1360 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG4 ( 1359 1346 )  100.n
R_D52103LOADxxQSG4 ( 0 1359 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG4 ( 1358 1346 )  100.n
R_D52104LOADxxQSG4 ( 0 1358 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG4 ( 1357 1346 )  100.n
R_D52105LOADxxQSG4 ( 0 1357 ) COMPLEX( 390., 0.)
R_D52107xxQSG4 ( 1356 1346 )  100.n
R_D52107LOADxxQSG4 ( 0 1356 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG4 ( 0 1355 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG4 ( 1355 1346 )  100.n
R_D52111xxQSG4 ( 1354 1346 )  100.n
R_D52111LOADxxQSG4 ( 1354 0 ) COMPLEX( 16.3926,-10.5885)
R_D52112xxQSG4 ( 1353 1346 )  100.n
R_D52112LOADxxQSG4 ( 1353 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG4 ( 1352 1346 )  100.n
R_D52113LOADxxQSG4 ( 1352 0 ) COMPLEX( 235.5726,-188.9955)
R_D52114xxQSG4 ( 1351 1346 )  100.n
R_D52114LOADxxQSG4 ( 1351 0 ) COMPLEX( 3.9963,-2.265)
R_D52115xxQSG4 ( 1350 1346 )  100.n
R_D52115LOADxxQSG4 ( 1350 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG4 ( 0 0 )  1.E+12
R_D52110xxQSG4 ( 1348 1346 )  100.n
R_D52110LOADxxQSG4 ( 1348 0 ) COMPLEX( 390., 0.)
R_D52109LOADxxQSG4 ( 0 1347 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG4 ( 1347 1346 )  100.n
R_D52106LOADxxQSG4 ( 1344 1345 )  100.n
R_D52106xxQSG4 ( 1345 1346 )  100.n
R_D52L2xxQSG4 ( 1303 1327 )  100.n
R_D52E2xxQSG4 ( 598 1327 )  100.n
R_D52E1xxQSG4 ( 614 1346 )  100.n
R_D52201xxQSG4 ( 1327 1342 )  100.n
R_D52201LOADxxQSG4 ( 0 1342 ) COMPLEX( 390., 0.)
R_D52202xxQSG4 ( 1341 1327 )  100.n
R_D52202LOADxxQSG4 ( 0 1341 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG4 ( 1340 1327 )  100.n
R_D52203LOADxxQSG4 ( 0 1340 ) COMPLEX( 123.9039,-92.928)
R_D52204xxQSG4 ( 1339 1327 )  100.n
R_D52204LOADxxQSG4 ( 0 1339 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG4 ( 1338 1327 )  100.n
R_D52205LOADxxQSG4 ( 0 1338 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG4 ( 1337 1327 )  100.n
R_D52206LOADxxQSG4 ( 1325 1337 )  100.n
R_D52208LOADxxQSG4 ( 0 1336 ) COMPLEX( 390., 0.)
R_D52208xxQSG4 ( 1336 1327 )  100.n
R_D52211xxQSG4 ( 1335 1327 )  100.n
R_D52211LOADxxQSG4 ( 1335 0 ) COMPLEX( 30.976, 0.)
R_D52212xxQSG4 ( 1334 1327 )  100.n
R_D52212LOADxxQSG4 ( 1334 0 ) COMPLEX( 390., 0.)
R_D52213xxQSG4 ( 1333 1327 )  100.n
R_D52213LOADxxQSG4 ( 1333 0 ) COMPLEX( 235.5726,-188.9955)
R_D52214xxQSG4 ( 1332 1327 )  100.n
R_D52214LOADxxQSG4 ( 1332 0 ) COMPLEX( 16.3926,-10.5885)
R_D52215xxQSG4 ( 1331 1327 )  100.n
R_D52215LOADxxQSG4 ( 1331 0 ) COMPLEX( 390., 0.)
R_D52216xxQSG4 ( 1330 1327 )  100.n
R_D52216LOADxxQSG4 ( 1330 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG4 ( 1329 1327 )  100.n
R_D52210LOADxxQSG4 ( 1329 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG4 ( 0 1328 ) COMPLEX( 390., 0.)
R_D52209xxQSG4 ( 1328 1327 )  100.n
R_D52207LOADxxQSG4 ( 1326 0 ) COMPLEX( 390., 0.)
R_D52207xxQSG4 ( 1326 1327 )  100.n
R_D52301xxQSG4 ( 1303 1324 )  100.n
R_D52301LOADxxQSG4 ( 0 1324 ) COMPLEX( 2.0445,-1.1034)
R_D52302xxQSG4 ( 1323 1303 )  100.n
R_D52302LOADxxQSG4 ( 0 1323 ) COMPLEX( 1.1652,-0.6288)
R_D52303xxQSG4 ( 1322 1303 )  100.n
R_D52303LOADxxQSG4 ( 0 1322 ) COMPLEX( 390., 0.)
R_D52304xxQSG4 ( 1321 1303 )  100.n
R_D52304LOADxxQSG4 ( 0 1321 ) COMPLEX( 1.7037,-0.9195)
R_D52305xxQSG4 ( 1320 1303 )  100.n
R_D52305LOADxxQSG4 ( 0 1320 ) COMPLEX( 390., 0.)
R_D52306xxQSG4 ( 1319 1303 )  100.n
R_D52306LOADxxQSG4 ( 0 1319 ) COMPLEX( 390., 0.)
R_D52308LOADxxQSG4 ( 0 1318 ) COMPLEX( 390., 0.)
R_D52308xxQSG4 ( 1318 1303 )  100.n
R_D52311xxQSG4 ( 1317 1303 )  100.n
R_D52311LOADxxQSG4 ( 1317 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG4 ( 1316 1303 )  100.n
R_D52312LOADxxQSG4 ( 1316 0 ) COMPLEX( 32.1234,-25.7721)
R_D52313xxQSG4 ( 1315 1303 )  100.n
R_D52313LOADxxQSG4 ( 1315 0 ) COMPLEX( 168.96,-126.72)
R_D52314xxQSG4 ( 1314 1303 )  100.n
R_D52314LOADxxQSG4 ( 1314 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG4 ( 1313 1303 )  100.n
R_D52315LOADxxQSG4 ( 1313 0 ) COMPLEX( 6.078,-3.2805)
R_D52316xxQSG4 ( 1312 1303 )  100.n
R_D52316LOADxxQSG4 ( 1312 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG4 ( 1311 1303 )  100.n
R_D52317LOADxxQSG4 ( 1311 0 ) COMPLEX( 4.2531,-2.5236)
R_D52310xxQSG4 ( 1310 1303 )  100.n
R_D52310LOADxxQSG4 ( 1310 0 ) COMPLEX( 2.4495,-0.8052)
R_D52318xxQSG4 ( 1309 1303 )  100.n
R_D52318LOADxxQSG4 ( 1309 0 ) COMPLEX( 2.2971,-1.3629)
R_D52319xxQSG4 ( 1308 1303 )  100.n
R_D52319LOADxxQSG4 ( 1308 0 ) COMPLEX( 20.4906,-13.2357)
R_D52309LOADxxQSG4 ( 0 1307 ) COMPLEX( 2.4495,-0.8052)
R_D52309xxQSG4 ( 1307 1303 )  100.n
R_D52307LOADxxQSG4 ( 1306 0 ) COMPLEX( 390., 0.)
R_D52307xxQSG4 ( 1306 1303 )  100.n
R_D52320xxQSG4 ( 1303 1305 )  100.n
R_D52320LOADxxQSG4 ( 0 1305 ) COMPLEX( 20.4906,-13.2357)
R_D52321xxQSG4 ( 1304 1303 )  100.n
R_D52321LOADxxQSG4 ( 0 1304 ) COMPLEX( 390., 0.)
R_D52322LOADxxQSG4 ( 0 1302 ) COMPLEX( 390., 0.)
R_D52322xxQSG4 ( 1302 1303 )  100.n
*-------------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U09CCM 
R_D52101xxU09 ( 1363 1395 )  100.n
R_D52101LOADxxU09 ( 0 1395 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU09 ( 1394 1363 )  100.n
R_D52102LOADxxU09 ( 0 1394 ) COMPLEX( 390., 0.)
R_D52103xxU09 ( 1393 1363 )  100.n
R_D52103LOADxxU09 ( 0 1393 ) COMPLEX( 390., 0.)
R_D52104xxU09 ( 1392 1363 )  100.n
R_D52104LOADxxU09 ( 0 1392 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU09 ( 1391 1363 )  100.n
R_D52105LOADxxU09 ( 0 1391 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU09 ( 1390 1363 )  100.n
R_D52106LOADxxU09 ( 0 1390 ) COMPLEX( 390., 0.)
R_D52107LOADxxU09 ( 0 1388 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU09 ( 0 1389 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU09 ( 1389 1363 )  100.n
R_D52107xxU09 ( 1388 1363 )  100.n
R_D52109xxU09 ( 1387 1363 )  100.n
R_D52109LOADxxU09 ( 1387 0 ) COMPLEX( 390., 0.)
R_D52110xxU09 ( 1386 1363 )  100.n
R_D52110LOADxxU09 ( 1386 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU09 ( 1385 1363 )  100.n
R_D52111LOADxxU09 ( 1385 0 ) COMPLEX( 390., 0.)
R_D52112xxU09 ( 1384 1363 )  100.n
R_D52112LOADxxU09 ( 1384 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU09 ( 1383 1363 )  100.n
R_D52113LOADxxU09 ( 1383 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU09 ( 1382 1363 )  100.n
R_D52114LOADxxU09 ( 1382 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU09 ( 1381 1363 )  100.n
R_D52116LOADxxU09 ( 1381 0 ) COMPLEX( 390., 0.)
R_D52ExxU09 ( 594 1363 )  100.n
R_D52115xxU09 ( 1379 1363 )  100.n
R_D52115LOADxxU09 ( 1379 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU09 ( 1363 1378 )  100.n
R_D52118LOADxxU09 ( 0 1378 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU09 ( 1377 1363 )  100.n
R_D52119LOADxxU09 ( 0 1377 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU09 ( 1376 1363 )  100.n
R_D52120LOADxxU09 ( 0 1376 ) COMPLEX( 390., 0.)
R_D52121xxU09 ( 1375 1363 )  100.n
R_D52121LOADxxU09 ( 0 1375 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU09 ( 1374 1363 )  100.n
R_D52122LOADxxU09 ( 0 1374 ) COMPLEX( 390., 0.)
R_D52123xxU09 ( 1373 1363 )  100.n
R_D52123LOADxxU09 ( 0 1373 ) COMPLEX( 390., 0.)
R_D52124LOADxxU09 ( 0 1371 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU09 ( 0 1372 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU09 ( 1372 1363 )  100.n
R_D52124xxU09 ( 1371 1363 )  100.n
R_D52125xxU09 ( 1370 1363 )  100.n
R_D52125LOADxxU09 ( 1370 0 ) COMPLEX( 390., 0.)
R_D52126xxU09 ( 1369 1363 )  100.n
R_D52126LOADxxU09 ( 1369 0 ) COMPLEX( 390., 0.)
R_D52127xxU09 ( 1368 1363 )  100.n
R_D52127LOADxxU09 ( 1368 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU09 ( 1367 1363 )  100.n
R_D52128LOADxxU09 ( 1367 0 ) COMPLEX( 390., 0.)
R_D52129xxU09 ( 1366 1363 )  100.n
R_D52129LOADxxU09 ( 1366 0 ) COMPLEX( 390., 0.)
R_D52130xxU09 ( 1365 1363 )  100.n
R_D52130LOADxxU09 ( 1365 0 ) COMPLEX( 390., 0.)
R_D52131xxU09 ( 1364 1363 )  100.n
R_D52131LOADxxU09 ( 1364 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU09 ( 1362 1363 )  100.n
R_D52132LOADxxU09 ( 1362 0 ) COMPLEX( 390., 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U10CCM 
R_D52101xxU10 ( 1397 1429 )  100.n
R_D52101LOADxxU10 ( 0 1429 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU10 ( 1428 1397 )  100.n
R_D52102LOADxxU10 ( 0 1428 ) COMPLEX( 390., 0.)
R_D52103xxU10 ( 1427 1397 )  100.n
R_D52103LOADxxU10 ( 0 1427 ) COMPLEX( 390., 0.)
R_D52104xxU10 ( 1426 1397 )  100.n
R_D52104LOADxxU10 ( 0 1426 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU10 ( 1425 1397 )  100.n
R_D52105LOADxxU10 ( 0 1425 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU10 ( 1424 1397 )  100.n
R_D52106LOADxxU10 ( 0 1424 ) COMPLEX( 390., 0.)
R_D52107LOADxxU10 ( 0 1422 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU10 ( 0 1423 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU10 ( 1423 1397 )  100.n
R_D52107xxU10 ( 1422 1397 )  100.n
R_D52109xxU10 ( 1421 1397 )  100.n
R_D52109LOADxxU10 ( 1421 0 ) COMPLEX( 390., 0.)
R_D52110xxU10 ( 1420 1397 )  100.n
R_D52110LOADxxU10 ( 1420 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU10 ( 1419 1397 )  100.n
R_D52111LOADxxU10 ( 1419 0 ) COMPLEX( 390., 0.)
R_D52112xxU10 ( 1418 1397 )  100.n
R_D52112LOADxxU10 ( 1418 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU10 ( 1417 1397 )  100.n
R_D52113LOADxxU10 ( 1417 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU10 ( 1416 1397 )  100.n
R_D52114LOADxxU10 ( 1416 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU10 ( 1415 1397 )  100.n
R_D52116LOADxxU10 ( 1415 0 ) COMPLEX( 390., 0.)
R_D52ExxU10 ( 596 1397 )  100.n
R_D52115xxU10 ( 1413 1397 )  100.n
R_D52115LOADxxU10 ( 1413 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU10 ( 1397 1412 )  100.n
R_D52118LOADxxU10 ( 0 1412 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU10 ( 1411 1397 )  100.n
R_D52119LOADxxU10 ( 0 1411 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU10 ( 1410 1397 )  100.n
R_D52120LOADxxU10 ( 0 1410 ) COMPLEX( 390., 0.)
R_D52121xxU10 ( 1409 1397 )  100.n
R_D52121LOADxxU10 ( 0 1409 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU10 ( 1408 1397 )  100.n
R_D52122LOADxxU10 ( 0 1408 ) COMPLEX( 390., 0.)
R_D52123xxU10 ( 1407 1397 )  100.n
R_D52123LOADxxU10 ( 0 1407 ) COMPLEX( 390., 0.)
R_D52124LOADxxU10 ( 0 1405 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU10 ( 0 1406 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU10 ( 1406 1397 )  100.n
R_D52124xxU10 ( 1405 1397 )  100.n
R_D52125xxU10 ( 1404 1397 )  100.n
R_D52125LOADxxU10 ( 1404 0 ) COMPLEX( 390., 0.)
R_D52126xxU10 ( 1403 1397 )  100.n
R_D52126LOADxxU10 ( 1403 0 ) COMPLEX( 390., 0.)
R_D52127xxU10 ( 1402 1397 )  100.n
R_D52127LOADxxU10 ( 1402 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU10 ( 1401 1397 )  100.n
R_D52128LOADxxU10 ( 1401 0 ) COMPLEX( 390., 0.)
R_D52129xxU10 ( 1400 1397 )  100.n
R_D52129LOADxxU10 ( 1400 0 ) COMPLEX( 390., 0.)
R_D52130xxU10 ( 1399 1397 )  100.n
R_D52130LOADxxU10 ( 1399 0 ) COMPLEX( 390., 0.)
R_D52131xxU10 ( 1398 1397 )  100.n
R_D52131LOADxxU10 ( 1398 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU10 ( 1396 1397 )  100.n
R_D52132LOADxxU10 ( 1396 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U11CCM 
R_D52101xxU11 ( 1431 1463 )  100.n
R_D52101LOADxxU11 ( 0 1463 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU11 ( 1462 1431 )  100.n
R_D52102LOADxxU11 ( 0 1462 ) COMPLEX( 390., 0.)
R_D52103xxU11 ( 1461 1431 )  100.n
R_D52103LOADxxU11 ( 0 1461 ) COMPLEX( 390., 0.)
R_D52104xxU11 ( 1460 1431 )  100.n
R_D52104LOADxxU11 ( 0 1460 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU11 ( 1459 1431 )  100.n
R_D52105LOADxxU11 ( 0 1459 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU11 ( 1458 1431 )  100.n
R_D52106LOADxxU11 ( 0 1458 ) COMPLEX( 390., 0.)
R_D52107LOADxxU11 ( 0 1456 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU11 ( 0 1457 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU11 ( 1457 1431 )  100.n
R_D52107xxU11 ( 1456 1431 )  100.n
R_D52109xxU11 ( 1455 1431 )  100.n
R_D52109LOADxxU11 ( 1455 0 ) COMPLEX( 390., 0.)
R_D52110xxU11 ( 1454 1431 )  100.n
R_D52110LOADxxU11 ( 1454 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU11 ( 1453 1431 )  100.n
R_D52111LOADxxU11 ( 1453 0 ) COMPLEX( 390., 0.)
R_D52112xxU11 ( 1452 1431 )  100.n
R_D52112LOADxxU11 ( 1452 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU11 ( 1451 1431 )  100.n
R_D52113LOADxxU11 ( 1451 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU11 ( 1450 1431 )  100.n
R_D52114LOADxxU11 ( 1450 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU11 ( 1449 1431 )  100.n
R_D52116LOADxxU11 ( 1449 0 ) COMPLEX( 390., 0.)
R_D52ExxU11 ( 600 1431 )  100.n
R_D52115xxU11 ( 1447 1431 )  100.n
R_D52115LOADxxU11 ( 1447 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU11 ( 1431 1446 )  100.n
R_D52118LOADxxU11 ( 0 1446 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU11 ( 1445 1431 )  100.n
R_D52119LOADxxU11 ( 0 1445 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU11 ( 1444 1431 )  100.n
R_D52120LOADxxU11 ( 0 1444 ) COMPLEX( 390., 0.)
R_D52121xxU11 ( 1443 1431 )  100.n
R_D52121LOADxxU11 ( 0 1443 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU11 ( 1442 1431 )  100.n
R_D52122LOADxxU11 ( 0 1442 ) COMPLEX( 390., 0.)
R_D52123xxU11 ( 1441 1431 )  100.n
R_D52123LOADxxU11 ( 0 1441 ) COMPLEX( 390., 0.)
R_D52124LOADxxU11 ( 0 1439 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU11 ( 0 1440 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU11 ( 1440 1431 )  100.n
R_D52124xxU11 ( 1439 1431 )  100.n
R_D52125xxU11 ( 1438 1431 )  100.n
R_D52125LOADxxU11 ( 1438 0 ) COMPLEX( 390., 0.)
R_D52126xxU11 ( 1437 1431 )  100.n
R_D52126LOADxxU11 ( 1437 0 ) COMPLEX( 390., 0.)
R_D52127xxU11 ( 1436 1431 )  100.n
R_D52127LOADxxU11 ( 1436 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU11 ( 1435 1431 )  100.n
R_D52128LOADxxU11 ( 1435 0 ) COMPLEX( 390., 0.)
R_D52129xxU11 ( 1434 1431 )  100.n
R_D52129LOADxxU11 ( 1434 0 ) COMPLEX( 390., 0.)
R_D52130xxU11 ( 1433 1431 )  100.n
R_D52130LOADxxU11 ( 1433 0 ) COMPLEX( 390., 0.)
R_D52131xxU11 ( 1432 1431 )  100.n
R_D52131LOADxxU11 ( 1432 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU11 ( 1430 1431 )  100.n
R_D52132LOADxxU11 ( 1430 0 ) COMPLEX( 390., 0.)
*---------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U12CCM 
R_D52101xxU12 ( 1465 1497 )  100.n
R_D52101LOADxxU12 ( 0 1497 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU12 ( 1496 1465 )  100.n
R_D52102LOADxxU12 ( 0 1496 ) COMPLEX( 390., 0.)
R_D52103xxU12 ( 1495 1465 )  100.n
R_D52103LOADxxU12 ( 0 1495 ) COMPLEX( 390., 0.)
R_D52104xxU12 ( 1494 1465 )  100.n
R_D52104LOADxxU12 ( 0 1494 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU12 ( 1493 1465 )  100.n
R_D52105LOADxxU12 ( 0 1493 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU12 ( 1492 1465 )  100.n
R_D52106LOADxxU12 ( 0 1492 ) COMPLEX( 390., 0.)
R_D52107LOADxxU12 ( 0 1490 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU12 ( 0 1491 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU12 ( 1491 1465 )  100.n
R_D52107xxU12 ( 1490 1465 )  100.n
R_D52109xxU12 ( 1489 1465 )  100.n
R_D52109LOADxxU12 ( 1489 0 ) COMPLEX( 390., 0.)
R_D52110xxU12 ( 1488 1465 )  100.n
R_D52110LOADxxU12 ( 1488 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU12 ( 1487 1465 )  100.n
R_D52111LOADxxU12 ( 1487 0 ) COMPLEX( 390., 0.)
R_D52112xxU12 ( 1486 1465 )  100.n
R_D52112LOADxxU12 ( 1486 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU12 ( 1485 1465 )  100.n
R_D52113LOADxxU12 ( 1485 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU12 ( 1484 1465 )  100.n
R_D52114LOADxxU12 ( 1484 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU12 ( 1483 1465 )  100.n
R_D52116LOADxxU12 ( 1483 0 ) COMPLEX( 390., 0.)
R_D52ExxU12 ( 599 1465 )  100.n
R_D52115xxU12 ( 1481 1465 )  100.n
R_D52115LOADxxU12 ( 1481 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU12 ( 1465 1480 )  100.n
R_D52118LOADxxU12 ( 0 1480 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU12 ( 1479 1465 )  100.n
R_D52119LOADxxU12 ( 0 1479 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU12 ( 1478 1465 )  100.n
R_D52120LOADxxU12 ( 0 1478 ) COMPLEX( 390., 0.)
R_D52121xxU12 ( 1477 1465 )  100.n
R_D52121LOADxxU12 ( 0 1477 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU12 ( 1476 1465 )  100.n
R_D52122LOADxxU12 ( 0 1476 ) COMPLEX( 390., 0.)
R_D52123xxU12 ( 1475 1465 )  100.n
R_D52123LOADxxU12 ( 0 1475 ) COMPLEX( 390., 0.)
R_D52124LOADxxU12 ( 0 1473 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU12 ( 0 1474 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU12 ( 1474 1465 )  100.n
R_D52124xxU12 ( 1473 1465 )  100.n
R_D52125xxU12 ( 1472 1465 )  100.n
R_D52125LOADxxU12 ( 1472 0 ) COMPLEX( 390., 0.)
R_D52126xxU12 ( 1471 1465 )  100.n
R_D52126LOADxxU12 ( 1471 0 ) COMPLEX( 390., 0.)
R_D52127xxU12 ( 1470 1465 )  100.n
R_D52127LOADxxU12 ( 1470 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU12 ( 1469 1465 )  100.n
R_D52128LOADxxU12 ( 1469 0 ) COMPLEX( 390., 0.)
R_D52129xxU12 ( 1468 1465 )  100.n
R_D52129LOADxxU12 ( 1468 0 ) COMPLEX( 390., 0.)
R_D52130xxU12 ( 1467 1465 )  100.n
R_D52130LOADxxU12 ( 1467 0 ) COMPLEX( 390., 0.)
R_D52131xxU12 ( 1466 1465 )  100.n
R_D52131LOADxxU12 ( 1466 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU12 ( 1464 1465 )  100.n
R_D52132LOADxxU12 ( 1464 0 ) COMPLEX( 390., 0.)
*------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA U13CCM 
R_D52101xxU13 ( 1499 1531 )  100.n
R_D52101LOADxxU13 ( 0 1531 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU13 ( 1530 1499 )  100.n
R_D52102LOADxxU13 ( 0 1530 ) COMPLEX( 390., 0.)
R_D52103xxU13 ( 1529 1499 )  100.n
R_D52103LOADxxU13 ( 0 1529 ) COMPLEX( 390., 0.)
R_D52104xxU13 ( 1528 1499 )  100.n
R_D52104LOADxxU13 ( 0 1528 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU13 ( 1527 1499 )  100.n
R_D52105LOADxxU13 ( 0 1527 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU13 ( 1526 1499 )  100.n
R_D52106LOADxxU13 ( 0 1526 ) COMPLEX( 390., 0.)
R_D52107LOADxxU13 ( 0 1524 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU13 ( 0 1525 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU13 ( 1525 1499 )  100.n
R_D52107xxU13 ( 1524 1499 )  100.n
R_D52109xxU13 ( 1523 1499 )  100.n
R_D52109LOADxxU13 ( 1523 0 ) COMPLEX( 390., 0.)
R_D52110xxU13 ( 1522 1499 )  100.n
R_D52110LOADxxU13 ( 1522 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU13 ( 1521 1499 )  100.n
R_D52111LOADxxU13 ( 1521 0 ) COMPLEX( 390., 0.)
R_D52112xxU13 ( 1520 1499 )  100.n
R_D52112LOADxxU13 ( 1520 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU13 ( 1519 1499 )  100.n
R_D52113LOADxxU13 ( 1519 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU13 ( 1518 1499 )  100.n
R_D52114LOADxxU13 ( 1518 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU13 ( 1517 1499 )  100.n
R_D52116LOADxxU13 ( 1517 0 ) COMPLEX( 390., 0.)
R_D52ExxU13 ( 617 1499 )  100.n
R_D52115xxU13 ( 1515 1499 )  100.n
R_D52115LOADxxU13 ( 1515 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU13 ( 1499 1514 )  100.n
R_D52118LOADxxU13 ( 0 1514 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU13 ( 1513 1499 )  100.n
R_D52119LOADxxU13 ( 0 1513 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU13 ( 1512 1499 )  100.n
R_D52120LOADxxU13 ( 0 1512 ) COMPLEX( 390., 0.)
R_D52121xxU13 ( 1511 1499 )  100.n
R_D52121LOADxxU13 ( 0 1511 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU13 ( 1510 1499 )  100.n
R_D52122LOADxxU13 ( 0 1510 ) COMPLEX( 390., 0.)
R_D52123xxU13 ( 1509 1499 )  100.n
R_D52123LOADxxU13 ( 0 1509 ) COMPLEX( 390., 0.)
R_D52124LOADxxU13 ( 0 1507 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU13 ( 0 1508 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU13 ( 1508 1499 )  100.n
R_D52124xxU13 ( 1507 1499 )  100.n
R_D52125xxU13 ( 1506 1499 )  100.n
R_D52125LOADxxU13 ( 1506 0 ) COMPLEX( 390., 0.)
R_D52126xxU13 ( 1505 1499 )  100.n
R_D52126LOADxxU13 ( 1505 0 ) COMPLEX( 390., 0.)
R_D52127xxU13 ( 1504 1499 )  100.n
R_D52127LOADxxU13 ( 1504 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU13 ( 1503 1499 )  100.n
R_D52128LOADxxU13 ( 1503 0 ) COMPLEX( 390., 0.)
R_D52129xxU13 ( 1502 1499 )  100.n
R_D52129LOADxxU13 ( 1502 0 ) COMPLEX( 390., 0.)
R_D52130xxU13 ( 1501 1499 )  100.n
R_D52130LOADxxU13 ( 1501 0 ) COMPLEX( 390., 0.)
R_D52131xxU13 ( 1500 1499 )  100.n
R_D52131LOADxxU13 ( 1500 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU13 ( 1498 1499 )  100.n
R_D52132LOADxxU13 ( 1498 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U14CCM 
R_D52101xxU14 ( 1533 1565 )  100.n
R_D52101LOADxxU14 ( 0 1565 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU14 ( 1564 1533 )  100.n
R_D52102LOADxxU14 ( 0 1564 ) COMPLEX( 390., 0.)
R_D52103xxU14 ( 1563 1533 )  100.n
R_D52103LOADxxU14 ( 0 1563 ) COMPLEX( 390., 0.)
R_D52104xxU14 ( 1562 1533 )  100.n
R_D52104LOADxxU14 ( 0 1562 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU14 ( 1561 1533 )  100.n
R_D52105LOADxxU14 ( 0 1561 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU14 ( 1560 1533 )  100.n
R_D52106LOADxxU14 ( 0 1560 ) COMPLEX( 390., 0.)
R_D52107LOADxxU14 ( 0 1558 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU14 ( 0 1559 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU14 ( 1559 1533 )  100.n
R_D52107xxU14 ( 1558 1533 )  100.n
R_D52109xxU14 ( 1557 1533 )  100.n
R_D52109LOADxxU14 ( 1557 0 ) COMPLEX( 390., 0.)
R_D52110xxU14 ( 1556 1533 )  100.n
R_D52110LOADxxU14 ( 1556 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU14 ( 1555 1533 )  100.n
R_D52111LOADxxU14 ( 1555 0 ) COMPLEX( 390., 0.)
R_D52112xxU14 ( 1554 1533 )  100.n
R_D52112LOADxxU14 ( 1554 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU14 ( 1553 1533 )  100.n
R_D52113LOADxxU14 ( 1553 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU14 ( 1552 1533 )  100.n
R_D52114LOADxxU14 ( 1552 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU14 ( 1551 1533 )  100.n
R_D52116LOADxxU14 ( 1551 0 ) COMPLEX( 390., 0.)
R_D52ExxU14 ( 615 1533 )  100.n
R_D52115xxU14 ( 1549 1533 )  100.n
R_D52115LOADxxU14 ( 1549 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU14 ( 1533 1548 )  100.n
R_D52118LOADxxU14 ( 0 1548 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU14 ( 1547 1533 )  100.n
R_D52119LOADxxU14 ( 0 1547 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU14 ( 1546 1533 )  100.n
R_D52120LOADxxU14 ( 0 1546 ) COMPLEX( 390., 0.)
R_D52121xxU14 ( 1545 1533 )  100.n
R_D52121LOADxxU14 ( 0 1545 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU14 ( 1544 1533 )  100.n
R_D52122LOADxxU14 ( 0 1544 ) COMPLEX( 390., 0.)
R_D52123xxU14 ( 1543 1533 )  100.n
R_D52123LOADxxU14 ( 0 1543 ) COMPLEX( 390., 0.)
R_D52124LOADxxU14 ( 0 1541 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU14 ( 0 1542 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU14 ( 1542 1533 )  100.n
R_D52124xxU14 ( 1541 1533 )  100.n
R_D52125xxU14 ( 1540 1533 )  100.n
R_D52125LOADxxU14 ( 1540 0 ) COMPLEX( 390., 0.)
R_D52126xxU14 ( 1539 1533 )  100.n
R_D52126LOADxxU14 ( 1539 0 ) COMPLEX( 390., 0.)
R_D52127xxU14 ( 1538 1533 )  100.n
R_D52127LOADxxU14 ( 1538 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU14 ( 1537 1533 )  100.n
R_D52128LOADxxU14 ( 1537 0 ) COMPLEX( 390., 0.)
R_D52129xxU14 ( 1536 1533 )  100.n
R_D52129LOADxxU14 ( 1536 0 ) COMPLEX( 390., 0.)
R_D52130xxU14 ( 1535 1533 )  100.n
R_D52130LOADxxU14 ( 1535 0 ) COMPLEX( 390., 0.)
R_D52131xxU14 ( 1534 1533 )  100.n
R_D52131LOADxxU14 ( 1534 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU14 ( 1532 1533 )  100.n
R_D52132LOADxxU14 ( 1532 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U15CCM 
R_D52101xxU15 ( 1567 1599 )  100.n
R_D52101LOADxxU15 ( 0 1599 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU15 ( 1598 1567 )  100.n
R_D52102LOADxxU15 ( 0 1598 ) COMPLEX( 390., 0.)
R_D52103xxU15 ( 1597 1567 )  100.n
R_D52103LOADxxU15 ( 0 1597 ) COMPLEX( 390., 0.)
R_D52104xxU15 ( 1596 1567 )  100.n
R_D52104LOADxxU15 ( 0 1596 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU15 ( 1595 1567 )  100.n
R_D52105LOADxxU15 ( 0 1595 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU15 ( 1594 1567 )  100.n
R_D52106LOADxxU15 ( 0 1594 ) COMPLEX( 390., 0.)
R_D52107LOADxxU15 ( 0 1592 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU15 ( 0 1593 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU15 ( 1593 1567 )  100.n
R_D52107xxU15 ( 1592 1567 )  100.n
R_D52109xxU15 ( 1591 1567 )  100.n
R_D52109LOADxxU15 ( 1591 0 ) COMPLEX( 390., 0.)
R_D52110xxU15 ( 1590 1567 )  100.n
R_D52110LOADxxU15 ( 1590 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU15 ( 1589 1567 )  100.n
R_D52111LOADxxU15 ( 1589 0 ) COMPLEX( 390., 0.)
R_D52112xxU15 ( 1588 1567 )  100.n
R_D52112LOADxxU15 ( 1588 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU15 ( 1587 1567 )  100.n
R_D52113LOADxxU15 ( 1587 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU15 ( 1586 1567 )  100.n
R_D52114LOADxxU15 ( 1586 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU15 ( 1585 1567 )  100.n
R_D52116LOADxxU15 ( 1585 0 ) COMPLEX( 390., 0.)
R_D52ExxU15 ( 621 1567 )  100.n
R_D52115xxU15 ( 1583 1567 )  100.n
R_D52115LOADxxU15 ( 1583 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU15 ( 1567 1582 )  100.n
R_D52118LOADxxU15 ( 0 1582 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU15 ( 1581 1567 )  100.n
R_D52119LOADxxU15 ( 0 1581 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU15 ( 1580 1567 )  100.n
R_D52120LOADxxU15 ( 0 1580 ) COMPLEX( 390., 0.)
R_D52121xxU15 ( 1579 1567 )  100.n
R_D52121LOADxxU15 ( 0 1579 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU15 ( 1578 1567 )  100.n
R_D52122LOADxxU15 ( 0 1578 ) COMPLEX( 390., 0.)
R_D52123xxU15 ( 1577 1567 )  100.n
R_D52123LOADxxU15 ( 0 1577 ) COMPLEX( 390., 0.)
R_D52124LOADxxU15 ( 0 1575 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU15 ( 0 1576 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU15 ( 1576 1567 )  100.n
R_D52124xxU15 ( 1575 1567 )  100.n
R_D52125xxU15 ( 1574 1567 )  100.n
R_D52125LOADxxU15 ( 1574 0 ) COMPLEX( 390., 0.)
R_D52126xxU15 ( 1573 1567 )  100.n
R_D52126LOADxxU15 ( 1573 0 ) COMPLEX( 390., 0.)
R_D52127xxU15 ( 1572 1567 )  100.n
R_D52127LOADxxU15 ( 1572 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU15 ( 1571 1567 )  100.n
R_D52128LOADxxU15 ( 1571 0 ) COMPLEX( 390., 0.)
R_D52129xxU15 ( 1570 1567 )  100.n
R_D52129LOADxxU15 ( 1570 0 ) COMPLEX( 390., 0.)
R_D52130xxU15 ( 1569 1567 )  100.n
R_D52130LOADxxU15 ( 1569 0 ) COMPLEX( 390., 0.)
R_D52131xxU15 ( 1568 1567 )  100.n
R_D52131LOADxxU15 ( 1568 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU15 ( 1566 1567 )  100.n
R_D52132LOADxxU15 ( 1566 0 ) COMPLEX( 390., 0.)
*------------------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA U16CCM 
R_D52101xxU16 ( 1601 1633 )  100.n
R_D52101LOADxxU16 ( 0 1633 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU16 ( 1632 1601 )  100.n
R_D52102LOADxxU16 ( 0 1632 ) COMPLEX( 390., 0.)
R_D52103xxU16 ( 1631 1601 )  100.n
R_D52103LOADxxU16 ( 0 1631 ) COMPLEX( 390., 0.)
R_D52104xxU16 ( 1630 1601 )  100.n
R_D52104LOADxxU16 ( 0 1630 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU16 ( 1629 1601 )  100.n
R_D52105LOADxxU16 ( 0 1629 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU16 ( 1628 1601 )  100.n
R_D52106LOADxxU16 ( 0 1628 ) COMPLEX( 390., 0.)
R_D52107LOADxxU16 ( 0 1626 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU16 ( 0 1627 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU16 ( 1627 1601 )  100.n
R_D52107xxU16 ( 1626 1601 )  100.n
R_D52109xxU16 ( 1625 1601 )  100.n
R_D52109LOADxxU16 ( 1625 0 ) COMPLEX( 390., 0.)
R_D52110xxU16 ( 1624 1601 )  100.n
R_D52110LOADxxU16 ( 1624 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU16 ( 1623 1601 )  100.n
R_D52111LOADxxU16 ( 1623 0 ) COMPLEX( 390., 0.)
R_D52112xxU16 ( 1622 1601 )  100.n
R_D52112LOADxxU16 ( 1622 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU16 ( 1621 1601 )  100.n
R_D52113LOADxxU16 ( 1621 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU16 ( 1620 1601 )  100.n
R_D52114LOADxxU16 ( 1620 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU16 ( 1619 1601 )  100.n
R_D52116LOADxxU16 ( 1619 0 ) COMPLEX( 390., 0.)
R_D52ExxU16 ( 620 1601 )  100.n
R_D52115xxU16 ( 1617 1601 )  100.n
R_D52115LOADxxU16 ( 1617 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU16 ( 1601 1616 )  100.n
R_D52118LOADxxU16 ( 0 1616 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU16 ( 1615 1601 )  100.n
R_D52119LOADxxU16 ( 0 1615 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU16 ( 1614 1601 )  100.n
R_D52120LOADxxU16 ( 0 1614 ) COMPLEX( 390., 0.)
R_D52121xxU16 ( 1613 1601 )  100.n
R_D52121LOADxxU16 ( 0 1613 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU16 ( 1612 1601 )  100.n
R_D52122LOADxxU16 ( 0 1612 ) COMPLEX( 390., 0.)
R_D52123xxU16 ( 1611 1601 )  100.n
R_D52123LOADxxU16 ( 0 1611 ) COMPLEX( 390., 0.)
R_D52124LOADxxU16 ( 0 1609 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU16 ( 0 1610 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU16 ( 1610 1601 )  100.n
R_D52124xxU16 ( 1609 1601 )  100.n
R_D52125xxU16 ( 1608 1601 )  100.n
R_D52125LOADxxU16 ( 1608 0 ) COMPLEX( 390., 0.)
R_D52126xxU16 ( 1607 1601 )  100.n
R_D52126LOADxxU16 ( 1607 0 ) COMPLEX( 390., 0.)
R_D52127xxU16 ( 1606 1601 )  100.n
R_D52127LOADxxU16 ( 1606 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU16 ( 1605 1601 )  100.n
R_D52128LOADxxU16 ( 1605 0 ) COMPLEX( 390., 0.)
R_D52129xxU16 ( 1604 1601 )  100.n
R_D52129LOADxxU16 ( 1604 0 ) COMPLEX( 390., 0.)
R_D52130xxU16 ( 1603 1601 )  100.n
R_D52130LOADxxU16 ( 1603 0 ) COMPLEX( 390., 0.)
R_D52131xxU16 ( 1602 1601 )  100.n
R_D52131LOADxxU16 ( 1602 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU16 ( 1600 1601 )  100.n
R_D52132LOADxxU16 ( 1600 0 ) COMPLEX( 390., 0.)
*------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSSE5 
R_D52L2xxQSSE5 ( 1634 1639 )  100.n
R_D52L1xxQSSE5 ( 0 0 )  1.E+12
R_D52101LOADxxQSSE5 ( 0 1635 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE5 ( 1635 1636 )  100.n
R_D52102LOADxxQSSE5 ( 0 1637 ) COMPLEX( 390., 0.)
R_D52102xxQSSE5 ( 1637 1636 )  100.n
R_D52201LOADxxQSSE5 ( 0 1638 ) COMPLEX( 9.7692,-5.5365)
R_D52201xxQSSE5 ( 1638 1639 )  100.n
R_D52202LOADxxQSSE5 ( 0 1640 ) COMPLEX( 390., 0.)
R_D52202xxQSSE5 ( 1640 1639 )  100.n
R_D52203LOADxxQSSE5 ( 0 1641 ) COMPLEX( 390., 0.)
R_D52203xxQSSE5 ( 1641 1639 )  100.n
R_D52301LOADxxQSSE5 ( 0 1642 ) COMPLEX( 10.7391,-6.372)
R_D52301xxQSSE5 ( 1642 1634 )  100.n
R_D52302LOADxxQSSE5 ( 0 1643 ) COMPLEX( 26.6742,-17.9253)
R_D52302xxQSSE5 ( 1643 1634 )  100.n
R_D52303LOADxxQSSE5 ( 0 1644 ) COMPLEX( 559.5039,-346.7493)
R_D52303xxQSSE5 ( 1644 1634 )  100.n
R_D52304LOADxxQSSE5 ( 0 1645 ) COMPLEX( 390., 0.)
R_D52304xxQSSE5 ( 1645 1634 )  100.n
R_D52305LOADxxQSSE5 ( 0 1646 ) COMPLEX( 390., 0.)
R_D52305xxQSSE5 ( 1646 1634 )  100.n
R_D52306LOADxxQSSE5 ( 0 1647 ) COMPLEX( 390., 0.)
R_D52306xxQSSE5 ( 1647 1634 )  100.n
R_D52E2xxQSSE5 ( 554 1639 )  100.n
R_D52E1xxQSSE5 ( 570 1636 )  100.n
*------------------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA QSSE6 
R_D52E1xxQSSE6 ( 558 1650 )  100.n
R_D52E2xxQSSE6 ( 578 1653 )  100.n
R_D52306xxQSSE6 ( 1661 1648 )  100.n
R_D52306LOADxxQSSE6 ( 0 1661 ) COMPLEX( 390., 0.)
R_D52305xxQSSE6 ( 1660 1648 )  100.n
R_D52305LOADxxQSSE6 ( 0 1660 ) COMPLEX( 390., 0.)
R_D52304xxQSSE6 ( 1659 1648 )  100.n
R_D52304LOADxxQSSE6 ( 0 1659 ) COMPLEX( 390., 0.)
R_D52303xxQSSE6 ( 1658 1648 )  100.n
R_D52303LOADxxQSSE6 ( 0 1658 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE6 ( 1657 1648 )  100.n
R_D52302LOADxxQSSE6 ( 0 1657 ) COMPLEX( 26.6742,-17.9253)
R_D52301xxQSSE6 ( 1656 1648 )  100.n
R_D52301LOADxxQSSE6 ( 0 1656 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE6 ( 1655 1653 )  100.n
R_D52203LOADxxQSSE6 ( 0 1655 ) COMPLEX( 390., 0.)
R_D52202xxQSSE6 ( 1654 1653 )  100.n
R_D52202LOADxxQSSE6 ( 0 1654 ) COMPLEX( 390., 0.)
R_D52201xxQSSE6 ( 1652 1653 )  100.n
R_D52201LOADxxQSSE6 ( 0 1652 ) COMPLEX( 9.7692,-5.5365)
R_D52102xxQSSE6 ( 1651 1650 )  100.n
R_D52102LOADxxQSSE6 ( 0 1651 ) COMPLEX( 390., 0.)
R_D52101xxQSSE6 ( 1649 1650 )  100.n
R_D52101LOADxxQSSE6 ( 0 1649 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE6 ( 0 0 )  1.E+12
R_D52L2xxQSSE6 ( 1648 1653 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSSE7 
R_D52E1xxQSSE7 ( 547 1664 )  100.n
R_D52E2xxQSSE7 ( 564 1668 )  100.n
R_D52307xxQSSE7 ( 1677 1662 )  100.n
R_D52307LOADxxQSSE7 ( 0 1677 ) COMPLEX( 13.9875,-8.6688)
R_D52306xxQSSE7 ( 1676 1662 )  100.n
R_D52306LOADxxQSSE7 ( 0 1676 ) COMPLEX( 390., 0.)
R_D52305xxQSSE7 ( 1675 1662 )  100.n
R_D52305LOADxxQSSE7 ( 0 1675 ) COMPLEX( 390., 0.)
R_D52304xxQSSE7 ( 1674 1662 )  100.n
R_D52304LOADxxQSSE7 ( 0 1674 ) COMPLEX( 390., 0.)
R_D52303xxQSSE7 ( 1673 1662 )  100.n
R_D52303LOADxxQSSE7 ( 0 1673 ) COMPLEX( 559.5039,-346.7493)
R_D52302xxQSSE7 ( 1672 1662 )  100.n
R_D52302LOADxxQSSE7 ( 0 1672 ) COMPLEX( 26.6742,-17.9253)
R_D52301xxQSSE7 ( 1671 1662 )  100.n
R_D52301LOADxxQSSE7 ( 0 1671 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE7 ( 1670 1668 )  100.n
R_D52203LOADxxQSSE7 ( 0 1670 ) COMPLEX( 390., 0.)
R_D52202xxQSSE7 ( 1669 1668 )  100.n
R_D52202LOADxxQSSE7 ( 0 1669 ) COMPLEX( 390., 0.)
R_D52201xxQSSE7 ( 1667 1668 )  100.n
R_D52201LOADxxQSSE7 ( 0 1667 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE7 ( 1666 1664 )  100.n
R_D52103LOADxxQSSE7 ( 0 1666 ) COMPLEX( 390., 0.)
R_D52102xxQSSE7 ( 1665 1664 )  100.n
R_D52102LOADxxQSSE7 ( 0 1665 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE7 ( 1663 1664 )  100.n
R_D52101LOADxxQSSE7 ( 0 1663 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE7 ( 0 0 )  1.E+12
R_D52L2xxQSSE7 ( 1662 1668 )  100.n
*------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSG5 
R_D52101xxQSG5 ( 1679 1740 )  100.n
R_D52101LOADxxQSG5 ( 0 1740 ) COMPLEX( 390., 0.)
R_D52102xxQSG5 ( 1739 1679 )  100.n
R_D52102LOADxxQSG5 ( 0 1739 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG5 ( 1738 1679 )  100.n
R_D52103LOADxxQSG5 ( 0 1738 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG5 ( 1737 1679 )  100.n
R_D52104LOADxxQSG5 ( 0 1737 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG5 ( 1736 1679 )  100.n
R_D52105LOADxxQSG5 ( 0 1736 ) COMPLEX( 390., 0.)
R_D52107xxQSG5 ( 1735 1679 )  100.n
R_D52107LOADxxQSG5 ( 0 1735 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG5 ( 0 1734 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG5 ( 1734 1679 )  100.n
R_D52111xxQSG5 ( 1733 1679 )  100.n
R_D52111LOADxxQSG5 ( 1733 0 ) COMPLEX( 16.3926,-10.5885)
R_D52112xxQSG5 ( 1732 1679 )  100.n
R_D52112LOADxxQSG5 ( 1732 0 ) COMPLEX( 235.5726,-188.9955)
R_D52113xxQSG5 ( 1731 1679 )  100.n
R_D52113LOADxxQSG5 ( 1731 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG5 ( 1730 1679 )  100.n
R_D52114LOADxxQSG5 ( 1730 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG5 ( 1729 1679 )  100.n
R_D52115LOADxxQSG5 ( 1729 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG5 ( 0 0 )  1.E+12
R_D52110xxQSG5 ( 1727 1679 )  100.n
R_D52110LOADxxQSG5 ( 1727 0 ) COMPLEX( 390., 0.)
R_D52109LOADxxQSG5 ( 0 1726 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG5 ( 1726 1679 )  100.n
R_D52106LOADxxQSG5 ( 1724 1725 )  100.n
R_D52106xxQSG5 ( 1725 1679 )  100.n
R_D52L2xxQSG5 ( 1681 1709 )  100.n
R_D52E2xxQSG5 ( 551 1709 )  100.n
R_D52E1xxQSG5 ( 569 1679 )  100.n
R_D52201xxQSG5 ( 1709 1722 )  100.n
R_D52201LOADxxQSG5 ( 0 1722 ) COMPLEX( 123.9039,-92.928)
R_D52202xxQSG5 ( 1721 1709 )  100.n
R_D52202LOADxxQSG5 ( 0 1721 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG5 ( 1720 1709 )  100.n
R_D52203LOADxxQSG5 ( 0 1720 ) COMPLEX( 390., 0.)
R_D52204xxQSG5 ( 1719 1709 )  100.n
R_D52204LOADxxQSG5 ( 0 1719 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG5 ( 1718 1709 )  100.n
R_D52205LOADxxQSG5 ( 0 1718 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG5 ( 1717 1709 )  100.n
R_D52206LOADxxQSG5 ( 1707 1717 )  100.n
R_D52208LOADxxQSG5 ( 0 1716 ) COMPLEX( 390., 0.)
R_D52208xxQSG5 ( 1716 1709 )  100.n
R_D52211xxQSG5 ( 1715 1709 )  100.n
R_D52211LOADxxQSG5 ( 1715 0 ) COMPLEX( 235.5726,-188.9955)
R_D52212xxQSG5 ( 1714 1709 )  100.n
R_D52212LOADxxQSG5 ( 1714 0 ) COMPLEX( 16.3926,-10.5885)
R_D52213xxQSG5 ( 1713 1709 )  100.n
R_D52213LOADxxQSG5 ( 1713 0 ) COMPLEX( 390., 0.)
R_D52214xxQSG5 ( 1712 1709 )  100.n
R_D52214LOADxxQSG5 ( 1712 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG5 ( 1711 1709 )  100.n
R_D52210LOADxxQSG5 ( 1711 0 ) COMPLEX( 30.976, 0.)
R_D52209LOADxxQSG5 ( 0 1710 ) COMPLEX( 390., 0.)
R_D52209xxQSG5 ( 1710 1709 )  100.n
R_D52207LOADxxQSG5 ( 1708 0 ) COMPLEX( 390., 0.)
R_D52207xxQSG5 ( 1708 1709 )  100.n
R_D52301xxQSG5 ( 1681 1706 )  100.n
R_D52301LOADxxQSG5 ( 0 1706 ) COMPLEX( 2.0445,-1.1034)
R_D52302xxQSG5 ( 1705 1681 )  100.n
R_D52302LOADxxQSG5 ( 0 1705 ) COMPLEX( 390., 0.)
R_D52303xxQSG5 ( 1704 1681 )  100.n
R_D52303LOADxxQSG5 ( 0 1704 ) COMPLEX( 176.6793,-141.7467)
R_D52304xxQSG5 ( 1703 1681 )  100.n
R_D52304LOADxxQSG5 ( 0 1703 ) COMPLEX( 390., 0.)
R_D52305xxQSG5 ( 1702 1681 )  100.n
R_D52305LOADxxQSG5 ( 0 1702 ) COMPLEX( 390., 0.)
R_D52306xxQSG5 ( 1701 1681 )  100.n
R_D52306LOADxxQSG5 ( 0 1701 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG5 ( 0 1700 ) COMPLEX( 390., 0.)
R_D52308xxQSG5 ( 1700 1681 )  100.n
R_D52311xxQSG5 ( 1699 1681 )  100.n
R_D52311LOADxxQSG5 ( 1699 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG5 ( 1698 1681 )  100.n
R_D52312LOADxxQSG5 ( 1698 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG5 ( 1697 1681 )  100.n
R_D52313LOADxxQSG5 ( 1697 0 ) COMPLEX( 168.96,-126.72)
R_D52314xxQSG5 ( 1696 1681 )  100.n
R_D52314LOADxxQSG5 ( 1696 0 ) COMPLEX( 168.96,-126.72)
R_D52315xxQSG5 ( 1695 1681 )  100.n
R_D52315LOADxxQSG5 ( 1695 0 ) COMPLEX( 390., 0.)
R_D52316xxQSG5 ( 1694 1681 )  100.n
R_D52316LOADxxQSG5 ( 1694 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG5 ( 1693 1681 )  100.n
R_D52317LOADxxQSG5 ( 1693 0 ) COMPLEX( 390., 0.)
R_D52310xxQSG5 ( 1692 1681 )  100.n
R_D52310LOADxxQSG5 ( 1692 0 ) COMPLEX( 390., 0.)
R_D52318xxQSG5 ( 1691 1681 )  100.n
R_D52318LOADxxQSG5 ( 1691 0 ) COMPLEX( 5.8614,-3.3219)
R_D52319xxQSG5 ( 1690 1681 )  100.n
R_D52319LOADxxQSG5 ( 1690 0 ) COMPLEX( 5.8614,-3.3219)
R_D52309LOADxxQSG5 ( 0 1689 ) COMPLEX( 390., 0.)
R_D52309xxQSG5 ( 1689 1681 )  100.n
R_D52307LOADxxQSG5 ( 1688 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG5 ( 1688 1681 )  100.n
R_D52320xxQSG5 ( 1681 1687 )  100.n
R_D52320LOADxxQSG5 ( 0 1687 ) COMPLEX( 390., 0.)
R_D52321xxQSG5 ( 1686 1681 )  100.n
R_D52321LOADxxQSG5 ( 0 1686 ) COMPLEX( 32.1234,-25.7721)
R_D52322LOADxxQSG5 ( 0 1685 ) COMPLEX( 32.1234,-25.7721)
R_D52322xxQSG5 ( 1685 1681 )  100.n
R_D52324xxQSG5 ( 1684 1681 )  100.n
R_D52324LOADxxQSG5 ( 1684 0 ) COMPLEX( 6.078,-3.2805)
R_D52325xxQSG5 ( 1683 1681 )  100.n
R_D52325LOADxxQSG5 ( 1683 0 ) COMPLEX( 20.4906,-13.2357)
R_D52326xxQSG5 ( 1682 1681 )  100.n
R_D52326LOADxxQSG5 ( 1682 0 ) COMPLEX( 20.4906,-13.2357)
R_D52323xxQSG5 ( 1680 1681 )  100.n
R_D52323LOADxxQSG5 ( 1680 0 ) COMPLEX( 6.078,-3.2805)
R_D52116xxQSG5 ( 1678 1679 )  100.n
R_D52116LOADxxQSG5 ( 1678 0 ) COMPLEX( 3.9963,-2.265)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSG6 
R_D52207xxQSG6 ( 1742 1743 )  100.n
R_D52207LOADxxQSG6 ( 1742 0 ) COMPLEX( 30.976, 0.)
R_D52209xxQSG6 ( 1744 1743 )  100.n
R_D52209LOADxxQSG6 ( 0 1744 ) COMPLEX( 390., 0.)
R_D52210LOADxxQSG6 ( 1745 0 ) COMPLEX( 390., 0.)
R_D52210xxQSG6 ( 1745 1743 )  100.n
R_D52215LOADxxQSG6 ( 1746 0 ) COMPLEX( 390., 0.)
R_D52215xxQSG6 ( 1746 1743 )  100.n
R_D52214LOADxxQSG6 ( 1747 0 ) COMPLEX( 16.3926,-10.5885)
R_D52214xxQSG6 ( 1747 1743 )  100.n
R_D52213LOADxxQSG6 ( 1748 0 ) COMPLEX( 235.5726,-188.9955)
R_D52213xxQSG6 ( 1748 1743 )  100.n
R_D52212LOADxxQSG6 ( 1749 0 ) COMPLEX( 235.5726,-188.9955)
R_D52212xxQSG6 ( 1749 1743 )  100.n
R_D52211LOADxxQSG6 ( 1750 0 ) COMPLEX( 235.5726,-188.9955)
R_D52211xxQSG6 ( 1750 1743 )  100.n
R_D52208xxQSG6 ( 1751 1743 )  100.n
R_D52208LOADxxQSG6 ( 0 1751 ) COMPLEX( 390., 0.)
R_D52206LOADxxQSG6 ( 1741 1752 )  100.n
R_D52206xxQSG6 ( 1752 1743 )  100.n
R_D52205LOADxxQSG6 ( 0 1753 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG6 ( 1753 1743 )  100.n
R_D52204LOADxxQSG6 ( 0 1754 ) COMPLEX( 3.9963,-2.265)
R_D52204xxQSG6 ( 1754 1743 )  100.n
R_D52203LOADxxQSG6 ( 0 1755 ) COMPLEX( 30.976, 0.)
R_D52203xxQSG6 ( 1755 1743 )  100.n
R_D52202LOADxxQSG6 ( 0 1756 ) COMPLEX( 86.7843,-60.576)
R_D52202xxQSG6 ( 1756 1743 )  100.n
R_D52201LOADxxQSG6 ( 0 1757 ) COMPLEX( 30.976, 0.)
R_D52201xxQSG6 ( 1743 1757 )  100.n
R_D52307xxQSG6 ( 1758 1759 )  100.n
R_D52307LOADxxQSG6 ( 1758 0 ) COMPLEX( 2.4495,-0.8052)
R_D52309xxQSG6 ( 1760 1759 )  100.n
R_D52309LOADxxQSG6 ( 0 1760 ) COMPLEX( 123.9039,-92.928)
R_D52310LOADxxQSG6 ( 1761 0 ) COMPLEX( 168.96,-126.72)
R_D52310xxQSG6 ( 1761 1759 )  100.n
R_D52317LOADxxQSG6 ( 1762 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG6 ( 1762 1759 )  100.n
R_D52316LOADxxQSG6 ( 1763 0 ) COMPLEX( 20.4906,-13.2357)
R_D52316xxQSG6 ( 1763 1759 )  100.n
R_D52315LOADxxQSG6 ( 1764 0 ) COMPLEX( 20.4906,-13.2357)
R_D52315xxQSG6 ( 1764 1759 )  100.n
R_D52314LOADxxQSG6 ( 1765 0 ) COMPLEX( 6.078,-3.2805)
R_D52314xxQSG6 ( 1765 1759 )  100.n
R_D52313LOADxxQSG6 ( 1766 0 ) COMPLEX( 6.078,-3.28)
R_D52313xxQSG6 ( 1766 1759 )  100.n
R_D52312LOADxxQSG6 ( 1767 0 ) COMPLEX( 64.2471,-51.5442)
R_D52312xxQSG6 ( 1767 1759 )  100.n
R_D52311LOADxxQSG6 ( 1768 0 ) COMPLEX( 390., 0.)
R_D52311xxQSG6 ( 1768 1759 )  100.n
R_D52308xxQSG6 ( 1769 1759 )  100.n
R_D52308LOADxxQSG6 ( 0 1769 ) COMPLEX( 390., 0.)
R_D52306LOADxxQSG6 ( 0 1770 ) COMPLEX( 2.4495,-0.8052)
R_D52306xxQSG6 ( 1770 1759 )  100.n
R_D52305LOADxxQSG6 ( 0 1771 ) COMPLEX( 390., 0.)
R_D52305xxQSG6 ( 1771 1759 )  100.n
R_D52304LOADxxQSG6 ( 0 1772 ) COMPLEX( 390., 0.)
R_D52304xxQSG6 ( 1772 1759 )  100.n
R_D52303LOADxxQSG6 ( 0 1773 ) COMPLEX( 6.078,-3.2805)
R_D52303xxQSG6 ( 1773 1759 )  100.n
R_D52302LOADxxQSG6 ( 0 1774 ) COMPLEX( 390., 0.)
R_D52302xxQSG6 ( 1774 1759 )  100.n
R_D52301LOADxxQSG6 ( 0 1775 ) COMPLEX( 2.0445,-1.1034)
R_D52301xxQSG6 ( 1759 1775 )  100.n
R_D52E1xxQSG6 ( 557 1779 )  100.n
R_D52E2xxQSG6 ( 574 1743 )  100.n
R_D52L2xxQSG6 ( 1759 1743 )  100.n
R_D52107xxQSG6 ( 1778 1779 )  100.n
R_D52107LOADxxQSG6 ( 1778 0 ) COMPLEX( 390., 0.)
R_D52109xxQSG6 ( 1780 1779 )  100.n
R_D52109LOADxxQSG6 ( 0 1780 ) COMPLEX( 3.9963,-2.265)
R_D52110LOADxxQSG6 ( 1781 0 ) COMPLEX( 390., 0.)
R_D52110xxQSG6 ( 1781 1779 )  100.n
R_D52L1xxQSG6 ( 0 0 )  1.E+12
R_D52113LOADxxQSG6 ( 1783 0 ) COMPLEX( 235.5726,-188.9955)
R_D52113xxQSG6 ( 1783 1779 )  100.n
R_D52112LOADxxQSG6 ( 1784 0 ) COMPLEX( 390., 0.)
R_D52112xxQSG6 ( 1784 1779 )  100.n
R_D52111LOADxxQSG6 ( 1785 0 ) COMPLEX( 16.3926,-10.5885)
R_D52111xxQSG6 ( 1785 1779 )  100.n
R_D52108xxQSG6 ( 1786 1779 )  100.n
R_D52108LOADxxQSG6 ( 0 1786 ) COMPLEX( 3.9963,-2.265)
R_D52106LOADxxQSG6 ( 1777 1787 )  100.n
R_D52106xxQSG6 ( 1787 1779 )  100.n
R_D52105LOADxxQSG6 ( 0 1788 ) COMPLEX( 390., 0.)
R_D52105xxQSG6 ( 1788 1779 )  100.n
R_D52104LOADxxQSG6 ( 0 1789 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG6 ( 1789 1779 )  100.n
R_D52103LOADxxQSG6 ( 0 1790 ) COMPLEX( 3.9963,-2.265)
R_D52103xxQSG6 ( 1790 1779 )  100.n
R_D52102LOADxxQSG6 ( 0 1791 ) COMPLEX( 86.7843,-60.576)
R_D52102xxQSG6 ( 1791 1779 )  100.n
R_D52101LOADxxQSG6 ( 0 1792 ) COMPLEX( 390., 0.)
R_D52101xxQSG6 ( 1779 1792 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSG7 
R_D52101xxQSG7 ( 1794 1860 )  100.n
R_D52101LOADxxQSG7 ( 0 1860 ) COMPLEX( 53.3484,-35.8503)
R_D52102xxQSG7 ( 1859 1794 )  100.n
R_D52102LOADxxQSG7 ( 0 1859 ) COMPLEX( 390., 0.)
R_D52103xxQSG7 ( 1858 1794 )  100.n
R_D52103LOADxxQSG7 ( 0 1858 ) COMPLEX( 86.7843,-60.576)
R_D52104xxQSG7 ( 1857 1794 )  100.n
R_D52104LOADxxQSG7 ( 0 1857 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG7 ( 1856 1794 )  100.n
R_D52105LOADxxQSG7 ( 0 1856 ) COMPLEX( 3.9963,-2.265)
R_D52106xxQSG7 ( 1855 1794 )  100.n
R_D52106LOADxxQSG7 ( 0 1855 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG7 ( 0 1854 ) COMPLEX( 390., 0.)
R_D52108xxQSG7 ( 1854 1794 )  100.n
R_D52112xxQSG7 ( 1853 1794 )  100.n
R_D52112LOADxxQSG7 ( 1853 0 ) COMPLEX( 102.99,-74.5635)
R_D52113xxQSG7 ( 1852 1794 )  100.n
R_D52113LOADxxQSG7 ( 1852 0 ) COMPLEX( 235.5726,-188.9955)
R_D52114xxQSG7 ( 1851 1794 )  100.n
R_D52114LOADxxQSG7 ( 1851 0 ) COMPLEX( 4.773,-2.832)
R_D52115xxQSG7 ( 1850 1794 )  100.n
R_D52115LOADxxQSG7 ( 1850 0 ) COMPLEX( 390., 0.)
R_D52116xxQSG7 ( 1849 1794 )  100.n
R_D52116LOADxxQSG7 ( 1849 0 ) COMPLEX( 390., 0.)
R_D52117xxQSG7 ( 1848 1794 )  100.n
R_D52117LOADxxQSG7 ( 1848 0 ) COMPLEX( 13.9875,-8.6688)
R_D52L1xxQSG7 ( 0 0 )  1.E+12
R_D52118xxQSG7 ( 1846 1794 )  100.n
R_D52118LOADxxQSG7 ( 1846 0 ) COMPLEX( 390., 0.)
R_D52111xxQSG7 ( 1845 1794 )  100.n
R_D52111LOADxxQSG7 ( 1845 0 ) COMPLEX( 390., 0.)
R_D52119xxQSG7 ( 1844 1794 )  100.n
R_D52119LOADxxQSG7 ( 1844 0 ) COMPLEX( 16.3926,-10.5885)
R_D52120xxQSG7 ( 1843 1794 )  100.n
R_D52120LOADxxQSG7 ( 1843 0 ) COMPLEX( 30.976, 0.)
R_D52109LOADxxQSG7 ( 0 1842 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG7 ( 1842 1794 )  100.n
R_D52107LOADxxQSG7 ( 1840 1841 )  100.n
R_D52107xxQSG7 ( 1841 1794 )  100.n
R_D52L2xxQSG7 ( 1796 1820 )  100.n
R_D52E2xxQSG7 ( 562 1820 )  100.n
R_D52E1xxQSG7 ( 546 1794 )  100.n
R_D52201xxQSG7 ( 1820 1838 )  100.n
R_D52201LOADxxQSG7 ( 0 1838 ) COMPLEX( 390., 0.)
R_D52202xxQSG7 ( 1837 1820 )  100.n
R_D52202LOADxxQSG7 ( 0 1837 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG7 ( 1836 1820 )  100.n
R_D52203LOADxxQSG7 ( 0 1836 ) COMPLEX( 123.9039,-92.928)
R_D52204xxQSG7 ( 1835 1820 )  100.n
R_D52204LOADxxQSG7 ( 0 1835 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG7 ( 1834 1820 )  100.n
R_D52205LOADxxQSG7 ( 0 1834 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG7 ( 1833 1820 )  100.n
R_D52206LOADxxQSG7 ( 1818 1833 )  100.n
R_D52208LOADxxQSG7 ( 0 1832 ) COMPLEX( 30.976, 0.)
R_D52208xxQSG7 ( 1832 1820 )  100.n
R_D52211xxQSG7 ( 1831 1820 )  100.n
R_D52211LOADxxQSG7 ( 1831 0 ) COMPLEX( 390., 0.)
R_D52212xxQSG7 ( 1830 1820 )  100.n
R_D52212LOADxxQSG7 ( 1830 0 ) COMPLEX( 390., 0.)
R_D52213xxQSG7 ( 1829 1820 )  100.n
R_D52213LOADxxQSG7 ( 1829 0 ) COMPLEX( 235.5726,-188.9955)
R_D52214xxQSG7 ( 1828 1820 )  100.n
R_D52214LOADxxQSG7 ( 1828 0 ) COMPLEX( 16.3926,-10.5885)
R_D52215xxQSG7 ( 1827 1820 )  100.n
R_D52215LOADxxQSG7 ( 1827 0 ) COMPLEX( 13.9875,-8.6688)
R_D52216xxQSG7 ( 1826 1820 )  100.n
R_D52216LOADxxQSG7 ( 1826 0 ) COMPLEX( 390., 0.)
R_D52217xxQSG7 ( 1825 1820 )  100.n
R_D52217LOADxxQSG7 ( 1825 0 ) COMPLEX( 390., 0.)
R_D52210xxQSG7 ( 1824 1820 )  100.n
R_D52210LOADxxQSG7 ( 1824 0 ) COMPLEX( 390., 0.)
R_D52218xxQSG7 ( 1823 1820 )  100.n
R_D52218LOADxxQSG7 ( 1823 0 ) COMPLEX( 30.976, 0.)
R_D52219xxQSG7 ( 1822 1820 )  100.n
R_D52219LOADxxQSG7 ( 1822 0 ) COMPLEX( 30.976, 0.)
R_D52209LOADxxQSG7 ( 0 1821 ) COMPLEX( 4.773,-2.832)
R_D52209xxQSG7 ( 1821 1820 )  100.n
R_D52207LOADxxQSG7 ( 1819 0 ) COMPLEX( 390., 0.)
R_D52207xxQSG7 ( 1819 1820 )  100.n
R_D52301xxQSG7 ( 1796 1817 )  100.n
R_D52301LOADxxQSG7 ( 0 1817 ) COMPLEX( 390., 0.)
R_D52302xxQSG7 ( 1816 1796 )  100.n
R_D52302LOADxxQSG7 ( 0 1816 ) COMPLEX( 176.6793,-141.7467)
R_D52303xxQSG7 ( 1815 1796 )  100.n
R_D52303LOADxxQSG7 ( 0 1815 ) COMPLEX( 390., 0.)
R_D52304xxQSG7 ( 1814 1796 )  100.n
R_D52304LOADxxQSG7 ( 0 1814 ) COMPLEX( 390., 0.)
R_D52305xxQSG7 ( 1813 1796 )  100.n
R_D52305LOADxxQSG7 ( 0 1813 ) COMPLEX( 2.4495,-0.8052)
R_D52306xxQSG7 ( 1812 1796 )  100.n
R_D52306LOADxxQSG7 ( 0 1812 ) COMPLEX( 390., 0.)
R_D52308LOADxxQSG7 ( 0 1811 ) COMPLEX( 390., 0.)
R_D52308xxQSG7 ( 1811 1796 )  100.n
R_D52311xxQSG7 ( 1810 1796 )  100.n
R_D52311LOADxxQSG7 ( 1810 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG7 ( 1809 1796 )  100.n
R_D52312LOADxxQSG7 ( 1809 0 ) COMPLEX( 390., 0.)
R_D52313xxQSG7 ( 1808 1796 )  100.n
R_D52313LOADxxQSG7 ( 1808 0 ) COMPLEX( 168.96,-126.72)
R_D52314xxQSG7 ( 1807 1796 )  100.n
R_D52314LOADxxQSG7 ( 1807 0 ) COMPLEX( 390., 0.)
R_D52315xxQSG7 ( 1806 1796 )  100.n
R_D52315LOADxxQSG7 ( 1806 0 ) COMPLEX( 2.4495,-0.8052)
R_D52316xxQSG7 ( 1805 1796 )  100.n
R_D52316LOADxxQSG7 ( 1805 0 ) COMPLEX( 64.2471,-51.5442)
R_D52317xxQSG7 ( 1804 1796 )  100.n
R_D52317LOADxxQSG7 ( 1804 0 ) COMPLEX( 6.078,-3.2805)
R_D52310xxQSG7 ( 1803 1796 )  100.n
R_D52310LOADxxQSG7 ( 1803 0 ) COMPLEX( 390., 0.)
R_D52318xxQSG7 ( 1802 1796 )  100.n
R_D52318LOADxxQSG7 ( 1802 0 ) COMPLEX( 6.078,-3.2805)
R_D52319xxQSG7 ( 1801 1796 )  100.n
R_D52319LOADxxQSG7 ( 1801 0 ) COMPLEX( 390., 0.)
R_D52309LOADxxQSG7 ( 0 1800 ) COMPLEX( 30.976, 0.)
R_D52309xxQSG7 ( 1800 1796 )  100.n
R_D52307LOADxxQSG7 ( 1799 0 ) COMPLEX( 390., 0.)
R_D52307xxQSG7 ( 1799 1796 )  100.n
R_D52320xxQSG7 ( 1796 1798 )  100.n
R_D52320LOADxxQSG7 ( 0 1798 ) COMPLEX( 20.4906,-13.2357)
R_D52321xxQSG7 ( 1797 1796 )  100.n
R_D52321LOADxxQSG7 ( 0 1797 ) COMPLEX( 20.4906,-13.2357)
R_D52322xxQSG7 ( 1795 1796 )  100.n
R_D52322LOADxxQSG7 ( 1795 0 ) COMPLEX( 390., 0.)
R_D52110LOADxxQSG7 ( 0 1793 ) COMPLEX( 3.9963,-2.265)
R_D52110xxQSG7 ( 1793 1794 )  100.n
*---------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U17CCM 
R_D52101xxU17 ( 1862 1894 )  100.n
R_D52101LOADxxU17 ( 0 1894 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU17 ( 1893 1862 )  100.n
R_D52102LOADxxU17 ( 0 1893 ) COMPLEX( 390., 0.)
R_D52103xxU17 ( 1892 1862 )  100.n
R_D52103LOADxxU17 ( 0 1892 ) COMPLEX( 390., 0.)
R_D52104xxU17 ( 1891 1862 )  100.n
R_D52104LOADxxU17 ( 0 1891 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU17 ( 1890 1862 )  100.n
R_D52105LOADxxU17 ( 0 1890 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU17 ( 1889 1862 )  100.n
R_D52106LOADxxU17 ( 0 1889 ) COMPLEX( 390., 0.)
R_D52107LOADxxU17 ( 0 1887 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU17 ( 0 1888 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU17 ( 1888 1862 )  100.n
R_D52107xxU17 ( 1887 1862 )  100.n
R_D52109xxU17 ( 1886 1862 )  100.n
R_D52109LOADxxU17 ( 1886 0 ) COMPLEX( 390., 0.)
R_D52110xxU17 ( 1885 1862 )  100.n
R_D52110LOADxxU17 ( 1885 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU17 ( 1884 1862 )  100.n
R_D52111LOADxxU17 ( 1884 0 ) COMPLEX( 390., 0.)
R_D52112xxU17 ( 1883 1862 )  100.n
R_D52112LOADxxU17 ( 1883 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU17 ( 1882 1862 )  100.n
R_D52113LOADxxU17 ( 1882 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU17 ( 1881 1862 )  100.n
R_D52114LOADxxU17 ( 1881 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU17 ( 1880 1862 )  100.n
R_D52116LOADxxU17 ( 1880 0 ) COMPLEX( 390., 0.)
R_D52ExxU17 ( 571 1862 )  100.n
R_D52115xxU17 ( 1878 1862 )  100.n
R_D52115LOADxxU17 ( 1878 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU17 ( 1862 1877 )  100.n
R_D52118LOADxxU17 ( 0 1877 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU17 ( 1876 1862 )  100.n
R_D52119LOADxxU17 ( 0 1876 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU17 ( 1875 1862 )  100.n
R_D52120LOADxxU17 ( 0 1875 ) COMPLEX( 390., 0.)
R_D52121xxU17 ( 1874 1862 )  100.n
R_D52121LOADxxU17 ( 0 1874 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU17 ( 1873 1862 )  100.n
R_D52122LOADxxU17 ( 0 1873 ) COMPLEX( 390., 0.)
R_D52123xxU17 ( 1872 1862 )  100.n
R_D52123LOADxxU17 ( 0 1872 ) COMPLEX( 390., 0.)
R_D52124LOADxxU17 ( 0 1870 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU17 ( 0 1871 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU17 ( 1871 1862 )  100.n
R_D52124xxU17 ( 1870 1862 )  100.n
R_D52125xxU17 ( 1869 1862 )  100.n
R_D52125LOADxxU17 ( 1869 0 ) COMPLEX( 390., 0.)
R_D52126xxU17 ( 1868 1862 )  100.n
R_D52126LOADxxU17 ( 1868 0 ) COMPLEX( 390., 0.)
R_D52127xxU17 ( 1867 1862 )  100.n
R_D52127LOADxxU17 ( 1867 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU17 ( 1866 1862 )  100.n
R_D52128LOADxxU17 ( 1866 0 ) COMPLEX( 390., 0.)
R_D52129xxU17 ( 1865 1862 )  100.n
R_D52129LOADxxU17 ( 1865 0 ) COMPLEX( 390., 0.)
R_D52130xxU17 ( 1864 1862 )  100.n
R_D52130LOADxxU17 ( 1864 0 ) COMPLEX( 390., 0.)
R_D52131xxU17 ( 1863 1862 )  100.n
R_D52131LOADxxU17 ( 1863 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU17 ( 1861 1862 )  100.n
R_D52132LOADxxU17 ( 1861 0 ) COMPLEX( 390., 0.)
*------------------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Aux CA U18CCM 
R_D52101xxU18 ( 1896 1928 )  100.n
R_D52101LOADxxU18 ( 0 1928 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU18 ( 1927 1896 )  100.n
R_D52102LOADxxU18 ( 0 1927 ) COMPLEX( 390., 0.)
R_D52103xxU18 ( 1926 1896 )  100.n
R_D52103LOADxxU18 ( 0 1926 ) COMPLEX( 390., 0.)
R_D52104xxU18 ( 1925 1896 )  100.n
R_D52104LOADxxU18 ( 0 1925 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU18 ( 1924 1896 )  100.n
R_D52105LOADxxU18 ( 0 1924 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU18 ( 1923 1896 )  100.n
R_D52106LOADxxU18 ( 0 1923 ) COMPLEX( 390., 0.)
R_D52107LOADxxU18 ( 0 1921 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU18 ( 0 1922 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU18 ( 1922 1896 )  100.n
R_D52107xxU18 ( 1921 1896 )  100.n
R_D52109xxU18 ( 1920 1896 )  100.n
R_D52109LOADxxU18 ( 1920 0 ) COMPLEX( 390., 0.)
R_D52110xxU18 ( 1919 1896 )  100.n
R_D52110LOADxxU18 ( 1919 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU18 ( 1918 1896 )  100.n
R_D52111LOADxxU18 ( 1918 0 ) COMPLEX( 390., 0.)
R_D52112xxU18 ( 1917 1896 )  100.n
R_D52112LOADxxU18 ( 1917 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU18 ( 1916 1896 )  100.n
R_D52113LOADxxU18 ( 1916 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU18 ( 1915 1896 )  100.n
R_D52114LOADxxU18 ( 1915 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU18 ( 1914 1896 )  100.n
R_D52116LOADxxU18 ( 1914 0 ) COMPLEX( 390., 0.)
R_D52ExxU18 ( 573 1896 )  100.n
R_D52115xxU18 ( 1912 1896 )  100.n
R_D52115LOADxxU18 ( 1912 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU18 ( 1896 1911 )  100.n
R_D52118LOADxxU18 ( 0 1911 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU18 ( 1910 1896 )  100.n
R_D52119LOADxxU18 ( 0 1910 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU18 ( 1909 1896 )  100.n
R_D52120LOADxxU18 ( 0 1909 ) COMPLEX( 390., 0.)
R_D52121xxU18 ( 1908 1896 )  100.n
R_D52121LOADxxU18 ( 0 1908 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU18 ( 1907 1896 )  100.n
R_D52122LOADxxU18 ( 0 1907 ) COMPLEX( 390., 0.)
R_D52123xxU18 ( 1906 1896 )  100.n
R_D52123LOADxxU18 ( 0 1906 ) COMPLEX( 390., 0.)
R_D52124LOADxxU18 ( 0 1904 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU18 ( 0 1905 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU18 ( 1905 1896 )  100.n
R_D52124xxU18 ( 1904 1896 )  100.n
R_D52125xxU18 ( 1903 1896 )  100.n
R_D52125LOADxxU18 ( 1903 0 ) COMPLEX( 390., 0.)
R_D52126xxU18 ( 1902 1896 )  100.n
R_D52126LOADxxU18 ( 1902 0 ) COMPLEX( 390., 0.)
R_D52127xxU18 ( 1901 1896 )  100.n
R_D52127LOADxxU18 ( 1901 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU18 ( 1900 1896 )  100.n
R_D52128LOADxxU18 ( 1900 0 ) COMPLEX( 390., 0.)
R_D52129xxU18 ( 1899 1896 )  100.n
R_D52129LOADxxU18 ( 1899 0 ) COMPLEX( 390., 0.)
R_D52130xxU18 ( 1898 1896 )  100.n
R_D52130LOADxxU18 ( 1898 0 ) COMPLEX( 390., 0.)
R_D52131xxU18 ( 1897 1896 )  100.n
R_D52131LOADxxU18 ( 1897 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU18 ( 1895 1896 )  100.n
R_D52132LOADxxU18 ( 1895 0 ) COMPLEX( 390., 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U19CCM 
R_D52101xxU19 ( 1930 1962 )  100.n
R_D52101LOADxxU19 ( 0 1962 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU19 ( 1961 1930 )  100.n
R_D52102LOADxxU19 ( 0 1961 ) COMPLEX( 390., 0.)
R_D52103xxU19 ( 1960 1930 )  100.n
R_D52103LOADxxU19 ( 0 1960 ) COMPLEX( 390., 0.)
R_D52104xxU19 ( 1959 1930 )  100.n
R_D52104LOADxxU19 ( 0 1959 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU19 ( 1958 1930 )  100.n
R_D52105LOADxxU19 ( 0 1958 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU19 ( 1957 1930 )  100.n
R_D52106LOADxxU19 ( 0 1957 ) COMPLEX( 390., 0.)
R_D52107LOADxxU19 ( 0 1955 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU19 ( 0 1956 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU19 ( 1956 1930 )  100.n
R_D52107xxU19 ( 1955 1930 )  100.n
R_D52109xxU19 ( 1954 1930 )  100.n
R_D52109LOADxxU19 ( 1954 0 ) COMPLEX( 390., 0.)
R_D52110xxU19 ( 1953 1930 )  100.n
R_D52110LOADxxU19 ( 1953 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU19 ( 1952 1930 )  100.n
R_D52111LOADxxU19 ( 1952 0 ) COMPLEX( 390., 0.)
R_D52112xxU19 ( 1951 1930 )  100.n
R_D52112LOADxxU19 ( 1951 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU19 ( 1950 1930 )  100.n
R_D52113LOADxxU19 ( 1950 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU19 ( 1949 1930 )  100.n
R_D52114LOADxxU19 ( 1949 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU19 ( 1948 1930 )  100.n
R_D52116LOADxxU19 ( 1948 0 ) COMPLEX( 390., 0.)
R_D52ExxU19 ( 577 1930 )  100.n
R_D52115xxU19 ( 1946 1930 )  100.n
R_D52115LOADxxU19 ( 1946 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU19 ( 1930 1945 )  100.n
R_D52118LOADxxU19 ( 0 1945 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU19 ( 1944 1930 )  100.n
R_D52119LOADxxU19 ( 0 1944 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU19 ( 1943 1930 )  100.n
R_D52120LOADxxU19 ( 0 1943 ) COMPLEX( 390., 0.)
R_D52121xxU19 ( 1942 1930 )  100.n
R_D52121LOADxxU19 ( 0 1942 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU19 ( 1941 1930 )  100.n
R_D52122LOADxxU19 ( 0 1941 ) COMPLEX( 390., 0.)
R_D52123xxU19 ( 1940 1930 )  100.n
R_D52123LOADxxU19 ( 0 1940 ) COMPLEX( 390., 0.)
R_D52124LOADxxU19 ( 0 1938 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU19 ( 0 1939 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU19 ( 1939 1930 )  100.n
R_D52124xxU19 ( 1938 1930 )  100.n
R_D52125xxU19 ( 1937 1930 )  100.n
R_D52125LOADxxU19 ( 1937 0 ) COMPLEX( 390., 0.)
R_D52126xxU19 ( 1936 1930 )  100.n
R_D52126LOADxxU19 ( 1936 0 ) COMPLEX( 390., 0.)
R_D52127xxU19 ( 1935 1930 )  100.n
R_D52127LOADxxU19 ( 1935 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU19 ( 1934 1930 )  100.n
R_D52128LOADxxU19 ( 1934 0 ) COMPLEX( 390., 0.)
R_D52129xxU19 ( 1933 1930 )  100.n
R_D52129LOADxxU19 ( 1933 0 ) COMPLEX( 390., 0.)
R_D52130xxU19 ( 1932 1930 )  100.n
R_D52130LOADxxU19 ( 1932 0 ) COMPLEX( 390., 0.)
R_D52131xxU19 ( 1931 1930 )  100.n
R_D52131LOADxxU19 ( 1931 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU19 ( 1929 1930 )  100.n
R_D52132LOADxxU19 ( 1929 0 ) COMPLEX( 390., 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U20CCM 
R_D52101xxU20 ( 1964 1996 )  100.n
R_D52101LOADxxU20 ( 0 1996 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU20 ( 1995 1964 )  100.n
R_D52102LOADxxU20 ( 0 1995 ) COMPLEX( 390., 0.)
R_D52103xxU20 ( 1994 1964 )  100.n
R_D52103LOADxxU20 ( 0 1994 ) COMPLEX( 390., 0.)
R_D52104xxU20 ( 1993 1964 )  100.n
R_D52104LOADxxU20 ( 0 1993 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU20 ( 1992 1964 )  100.n
R_D52105LOADxxU20 ( 0 1992 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU20 ( 1991 1964 )  100.n
R_D52106LOADxxU20 ( 0 1991 ) COMPLEX( 390., 0.)
R_D52107LOADxxU20 ( 0 1989 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU20 ( 0 1990 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU20 ( 1990 1964 )  100.n
R_D52107xxU20 ( 1989 1964 )  100.n
R_D52109xxU20 ( 1988 1964 )  100.n
R_D52109LOADxxU20 ( 1988 0 ) COMPLEX( 390., 0.)
R_D52110xxU20 ( 1987 1964 )  100.n
R_D52110LOADxxU20 ( 1987 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU20 ( 1986 1964 )  100.n
R_D52111LOADxxU20 ( 1986 0 ) COMPLEX( 390., 0.)
R_D52112xxU20 ( 1985 1964 )  100.n
R_D52112LOADxxU20 ( 1985 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU20 ( 1984 1964 )  100.n
R_D52113LOADxxU20 ( 1984 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU20 ( 1983 1964 )  100.n
R_D52114LOADxxU20 ( 1983 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU20 ( 1982 1964 )  100.n
R_D52116LOADxxU20 ( 1982 0 ) COMPLEX( 390., 0.)
R_D52ExxU20 ( 576 1964 )  100.n
R_D52115xxU20 ( 1980 1964 )  100.n
R_D52115LOADxxU20 ( 1980 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU20 ( 1964 1979 )  100.n
R_D52118LOADxxU20 ( 0 1979 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU20 ( 1978 1964 )  100.n
R_D52119LOADxxU20 ( 0 1978 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU20 ( 1977 1964 )  100.n
R_D52120LOADxxU20 ( 0 1977 ) COMPLEX( 390., 0.)
R_D52121xxU20 ( 1976 1964 )  100.n
R_D52121LOADxxU20 ( 0 1976 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU20 ( 1975 1964 )  100.n
R_D52122LOADxxU20 ( 0 1975 ) COMPLEX( 390., 0.)
R_D52123xxU20 ( 1974 1964 )  100.n
R_D52123LOADxxU20 ( 0 1974 ) COMPLEX( 390., 0.)
R_D52124LOADxxU20 ( 0 1972 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU20 ( 0 1973 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU20 ( 1973 1964 )  100.n
R_D52124xxU20 ( 1972 1964 )  100.n
R_D52125xxU20 ( 1971 1964 )  100.n
R_D52125LOADxxU20 ( 1971 0 ) COMPLEX( 390., 0.)
R_D52126xxU20 ( 1970 1964 )  100.n
R_D52126LOADxxU20 ( 1970 0 ) COMPLEX( 390., 0.)
R_D52127xxU20 ( 1969 1964 )  100.n
R_D52127LOADxxU20 ( 1969 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU20 ( 1968 1964 )  100.n
R_D52128LOADxxU20 ( 1968 0 ) COMPLEX( 390., 0.)
R_D52129xxU20 ( 1967 1964 )  100.n
R_D52129LOADxxU20 ( 1967 0 ) COMPLEX( 390., 0.)
R_D52130xxU20 ( 1966 1964 )  100.n
R_D52130LOADxxU20 ( 1966 0 ) COMPLEX( 390., 0.)
R_D52131xxU20 ( 1965 1964 )  100.n
R_D52131LOADxxU20 ( 1965 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU20 ( 1963 1964 )  100.n
R_D52132LOADxxU20 ( 1963 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U21CCM 
R_D52101xxU21 ( 1998 2030 )  100.n
R_D52101LOADxxU21 ( 0 2030 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU21 ( 2029 1998 )  100.n
R_D52102LOADxxU21 ( 0 2029 ) COMPLEX( 390., 0.)
R_D52103xxU21 ( 2028 1998 )  100.n
R_D52103LOADxxU21 ( 0 2028 ) COMPLEX( 390., 0.)
R_D52104xxU21 ( 2027 1998 )  100.n
R_D52104LOADxxU21 ( 0 2027 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU21 ( 2026 1998 )  100.n
R_D52105LOADxxU21 ( 0 2026 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU21 ( 2025 1998 )  100.n
R_D52106LOADxxU21 ( 0 2025 ) COMPLEX( 390., 0.)
R_D52107LOADxxU21 ( 0 2023 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU21 ( 0 2024 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU21 ( 2024 1998 )  100.n
R_D52107xxU21 ( 2023 1998 )  100.n
R_D52109xxU21 ( 2022 1998 )  100.n
R_D52109LOADxxU21 ( 2022 0 ) COMPLEX( 390., 0.)
R_D52110xxU21 ( 2021 1998 )  100.n
R_D52110LOADxxU21 ( 2021 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU21 ( 2020 1998 )  100.n
R_D52111LOADxxU21 ( 2020 0 ) COMPLEX( 390., 0.)
R_D52112xxU21 ( 2019 1998 )  100.n
R_D52112LOADxxU21 ( 2019 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU21 ( 2018 1998 )  100.n
R_D52113LOADxxU21 ( 2018 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU21 ( 2017 1998 )  100.n
R_D52114LOADxxU21 ( 2017 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU21 ( 2016 1998 )  100.n
R_D52116LOADxxU21 ( 2016 0 ) COMPLEX( 390., 0.)
R_D52ExxU21 ( 559 1998 )  100.n
R_D52115xxU21 ( 2014 1998 )  100.n
R_D52115LOADxxU21 ( 2014 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU21 ( 1998 2013 )  100.n
R_D52118LOADxxU21 ( 0 2013 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU21 ( 2012 1998 )  100.n
R_D52119LOADxxU21 ( 0 2012 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU21 ( 2011 1998 )  100.n
R_D52120LOADxxU21 ( 0 2011 ) COMPLEX( 390., 0.)
R_D52121xxU21 ( 2010 1998 )  100.n
R_D52121LOADxxU21 ( 0 2010 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU21 ( 2009 1998 )  100.n
R_D52122LOADxxU21 ( 0 2009 ) COMPLEX( 390., 0.)
R_D52123xxU21 ( 2008 1998 )  100.n
R_D52123LOADxxU21 ( 0 2008 ) COMPLEX( 390., 0.)
R_D52124LOADxxU21 ( 0 2006 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU21 ( 0 2007 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU21 ( 2007 1998 )  100.n
R_D52124xxU21 ( 2006 1998 )  100.n
R_D52125xxU21 ( 2005 1998 )  100.n
R_D52125LOADxxU21 ( 2005 0 ) COMPLEX( 390., 0.)
R_D52126xxU21 ( 2004 1998 )  100.n
R_D52126LOADxxU21 ( 2004 0 ) COMPLEX( 390., 0.)
R_D52127xxU21 ( 2003 1998 )  100.n
R_D52127LOADxxU21 ( 2003 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU21 ( 2002 1998 )  100.n
R_D52128LOADxxU21 ( 2002 0 ) COMPLEX( 390., 0.)
R_D52129xxU21 ( 2001 1998 )  100.n
R_D52129LOADxxU21 ( 2001 0 ) COMPLEX( 390., 0.)
R_D52130xxU21 ( 2000 1998 )  100.n
R_D52130LOADxxU21 ( 2000 0 ) COMPLEX( 390., 0.)
R_D52131xxU21 ( 1999 1998 )  100.n
R_D52131LOADxxU21 ( 1999 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU21 ( 1997 1998 )  100.n
R_D52132LOADxxU21 ( 1997 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U22CCM 
R_D52101xxU22 ( 2032 2064 )  100.n
R_D52101LOADxxU22 ( 0 2064 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU22 ( 2063 2032 )  100.n
R_D52102LOADxxU22 ( 0 2063 ) COMPLEX( 390., 0.)
R_D52103xxU22 ( 2062 2032 )  100.n
R_D52103LOADxxU22 ( 0 2062 ) COMPLEX( 390., 0.)
R_D52104xxU22 ( 2061 2032 )  100.n
R_D52104LOADxxU22 ( 0 2061 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU22 ( 2060 2032 )  100.n
R_D52105LOADxxU22 ( 0 2060 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU22 ( 2059 2032 )  100.n
R_D52106LOADxxU22 ( 0 2059 ) COMPLEX( 390., 0.)
R_D52107LOADxxU22 ( 0 2057 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU22 ( 0 2058 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU22 ( 2058 2032 )  100.n
R_D52107xxU22 ( 2057 2032 )  100.n
R_D52109xxU22 ( 2056 2032 )  100.n
R_D52109LOADxxU22 ( 2056 0 ) COMPLEX( 390., 0.)
R_D52110xxU22 ( 2055 2032 )  100.n
R_D52110LOADxxU22 ( 2055 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU22 ( 2054 2032 )  100.n
R_D52111LOADxxU22 ( 2054 0 ) COMPLEX( 390., 0.)
R_D52112xxU22 ( 2053 2032 )  100.n
R_D52112LOADxxU22 ( 2053 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU22 ( 2052 2032 )  100.n
R_D52113LOADxxU22 ( 2052 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU22 ( 2051 2032 )  100.n
R_D52114LOADxxU22 ( 2051 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU22 ( 2050 2032 )  100.n
R_D52116LOADxxU22 ( 2050 0 ) COMPLEX( 390., 0.)
R_D52ExxU22 ( 561 2032 )  100.n
R_D52115xxU22 ( 2048 2032 )  100.n
R_D52115LOADxxU22 ( 2048 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU22 ( 2032 2047 )  100.n
R_D52118LOADxxU22 ( 0 2047 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU22 ( 2046 2032 )  100.n
R_D52119LOADxxU22 ( 0 2046 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU22 ( 2045 2032 )  100.n
R_D52120LOADxxU22 ( 0 2045 ) COMPLEX( 390., 0.)
R_D52121xxU22 ( 2044 2032 )  100.n
R_D52121LOADxxU22 ( 0 2044 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU22 ( 2043 2032 )  100.n
R_D52122LOADxxU22 ( 0 2043 ) COMPLEX( 390., 0.)
R_D52123xxU22 ( 2042 2032 )  100.n
R_D52123LOADxxU22 ( 0 2042 ) COMPLEX( 390., 0.)
R_D52124LOADxxU22 ( 0 2040 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU22 ( 0 2041 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU22 ( 2041 2032 )  100.n
R_D52124xxU22 ( 2040 2032 )  100.n
R_D52125xxU22 ( 2039 2032 )  100.n
R_D52125LOADxxU22 ( 2039 0 ) COMPLEX( 390., 0.)
R_D52126xxU22 ( 2038 2032 )  100.n
R_D52126LOADxxU22 ( 2038 0 ) COMPLEX( 390., 0.)
R_D52127xxU22 ( 2037 2032 )  100.n
R_D52127LOADxxU22 ( 2037 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU22 ( 2036 2032 )  100.n
R_D52128LOADxxU22 ( 2036 0 ) COMPLEX( 390., 0.)
R_D52129xxU22 ( 2035 2032 )  100.n
R_D52129LOADxxU22 ( 2035 0 ) COMPLEX( 390., 0.)
R_D52130xxU22 ( 2034 2032 )  100.n
R_D52130LOADxxU22 ( 2034 0 ) COMPLEX( 390., 0.)
R_D52131xxU22 ( 2033 2032 )  100.n
R_D52131LOADxxU22 ( 2033 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU22 ( 2031 2032 )  100.n
R_D52132LOADxxU22 ( 2031 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U23CCM 
R_D52101xxU23 ( 2066 2098 )  100.n
R_D52101LOADxxU23 ( 0 2098 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU23 ( 2097 2066 )  100.n
R_D52102LOADxxU23 ( 0 2097 ) COMPLEX( 390., 0.)
R_D52103xxU23 ( 2096 2066 )  100.n
R_D52103LOADxxU23 ( 0 2096 ) COMPLEX( 390., 0.)
R_D52104xxU23 ( 2095 2066 )  100.n
R_D52104LOADxxU23 ( 0 2095 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU23 ( 2094 2066 )  100.n
R_D52105LOADxxU23 ( 0 2094 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU23 ( 2093 2066 )  100.n
R_D52106LOADxxU23 ( 0 2093 ) COMPLEX( 390., 0.)
R_D52107LOADxxU23 ( 0 2091 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU23 ( 0 2092 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU23 ( 2092 2066 )  100.n
R_D52107xxU23 ( 2091 2066 )  100.n
R_D52109xxU23 ( 2090 2066 )  100.n
R_D52109LOADxxU23 ( 2090 0 ) COMPLEX( 390., 0.)
R_D52110xxU23 ( 2089 2066 )  100.n
R_D52110LOADxxU23 ( 2089 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU23 ( 2088 2066 )  100.n
R_D52111LOADxxU23 ( 2088 0 ) COMPLEX( 390., 0.)
R_D52112xxU23 ( 2087 2066 )  100.n
R_D52112LOADxxU23 ( 2087 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU23 ( 2086 2066 )  100.n
R_D52113LOADxxU23 ( 2086 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU23 ( 2085 2066 )  100.n
R_D52114LOADxxU23 ( 2085 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU23 ( 2084 2066 )  100.n
R_D52116LOADxxU23 ( 2084 0 ) COMPLEX( 390., 0.)
R_D52ExxU23 ( 566 2066 )  100.n
R_D52115xxU23 ( 2082 2066 )  100.n
R_D52115LOADxxU23 ( 2082 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU23 ( 2066 2081 )  100.n
R_D52118LOADxxU23 ( 0 2081 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU23 ( 2080 2066 )  100.n
R_D52119LOADxxU23 ( 0 2080 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU23 ( 2079 2066 )  100.n
R_D52120LOADxxU23 ( 0 2079 ) COMPLEX( 390., 0.)
R_D52121xxU23 ( 2078 2066 )  100.n
R_D52121LOADxxU23 ( 0 2078 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU23 ( 2077 2066 )  100.n
R_D52122LOADxxU23 ( 0 2077 ) COMPLEX( 390., 0.)
R_D52123xxU23 ( 2076 2066 )  100.n
R_D52123LOADxxU23 ( 0 2076 ) COMPLEX( 390., 0.)
R_D52124LOADxxU23 ( 0 2074 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU23 ( 0 2075 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU23 ( 2075 2066 )  100.n
R_D52124xxU23 ( 2074 2066 )  100.n
R_D52125xxU23 ( 2073 2066 )  100.n
R_D52125LOADxxU23 ( 2073 0 ) COMPLEX( 390., 0.)
R_D52126xxU23 ( 2072 2066 )  100.n
R_D52126LOADxxU23 ( 2072 0 ) COMPLEX( 390., 0.)
R_D52127xxU23 ( 2071 2066 )  100.n
R_D52127LOADxxU23 ( 2071 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU23 ( 2070 2066 )  100.n
R_D52128LOADxxU23 ( 2070 0 ) COMPLEX( 390., 0.)
R_D52129xxU23 ( 2069 2066 )  100.n
R_D52129LOADxxU23 ( 2069 0 ) COMPLEX( 390., 0.)
R_D52130xxU23 ( 2068 2066 )  100.n
R_D52130LOADxxU23 ( 2068 0 ) COMPLEX( 390., 0.)
R_D52131xxU23 ( 2067 2066 )  100.n
R_D52131LOADxxU23 ( 2067 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU23 ( 2065 2066 )  100.n
R_D52132LOADxxU23 ( 2065 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U24CCM 
R_D52101xxU24 ( 2100 2132 )  100.n
R_D52101LOADxxU24 ( 0 2132 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU24 ( 2131 2100 )  100.n
R_D52102LOADxxU24 ( 0 2131 ) COMPLEX( 390., 0.)
R_D52103xxU24 ( 2130 2100 )  100.n
R_D52103LOADxxU24 ( 0 2130 ) COMPLEX( 390., 0.)
R_D52104xxU24 ( 2129 2100 )  100.n
R_D52104LOADxxU24 ( 0 2129 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU24 ( 2128 2100 )  100.n
R_D52105LOADxxU24 ( 0 2128 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU24 ( 2127 2100 )  100.n
R_D52106LOADxxU24 ( 0 2127 ) COMPLEX( 390., 0.)
R_D52107LOADxxU24 ( 0 2125 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU24 ( 0 2126 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU24 ( 2126 2100 )  100.n
R_D52107xxU24 ( 2125 2100 )  100.n
R_D52109xxU24 ( 2124 2100 )  100.n
R_D52109LOADxxU24 ( 2124 0 ) COMPLEX( 390., 0.)
R_D52110xxU24 ( 2123 2100 )  100.n
R_D52110LOADxxU24 ( 2123 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU24 ( 2122 2100 )  100.n
R_D52111LOADxxU24 ( 2122 0 ) COMPLEX( 390., 0.)
R_D52112xxU24 ( 2121 2100 )  100.n
R_D52112LOADxxU24 ( 2121 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU24 ( 2120 2100 )  100.n
R_D52113LOADxxU24 ( 2120 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU24 ( 2119 2100 )  100.n
R_D52114LOADxxU24 ( 2119 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU24 ( 2118 2100 )  100.n
R_D52116LOADxxU24 ( 2118 0 ) COMPLEX( 390., 0.)
R_D52ExxU24 ( 555 2100 )  100.n
R_D52115xxU24 ( 2116 2100 )  100.n
R_D52115LOADxxU24 ( 2116 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU24 ( 2100 2115 )  100.n
R_D52118LOADxxU24 ( 0 2115 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU24 ( 2114 2100 )  100.n
R_D52119LOADxxU24 ( 0 2114 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU24 ( 2113 2100 )  100.n
R_D52120LOADxxU24 ( 0 2113 ) COMPLEX( 390., 0.)
R_D52121xxU24 ( 2112 2100 )  100.n
R_D52121LOADxxU24 ( 0 2112 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU24 ( 2111 2100 )  100.n
R_D52122LOADxxU24 ( 0 2111 ) COMPLEX( 390., 0.)
R_D52123xxU24 ( 2110 2100 )  100.n
R_D52123LOADxxU24 ( 0 2110 ) COMPLEX( 390., 0.)
R_D52124LOADxxU24 ( 0 2108 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU24 ( 0 2109 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU24 ( 2109 2100 )  100.n
R_D52124xxU24 ( 2108 2100 )  100.n
R_D52125xxU24 ( 2107 2100 )  100.n
R_D52125LOADxxU24 ( 2107 0 ) COMPLEX( 390., 0.)
R_D52126xxU24 ( 2106 2100 )  100.n
R_D52126LOADxxU24 ( 2106 0 ) COMPLEX( 390., 0.)
R_D52127xxU24 ( 2105 2100 )  100.n
R_D52127LOADxxU24 ( 2105 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU24 ( 2104 2100 )  100.n
R_D52128LOADxxU24 ( 2104 0 ) COMPLEX( 390., 0.)
R_D52129xxU24 ( 2103 2100 )  100.n
R_D52129LOADxxU24 ( 2103 0 ) COMPLEX( 390., 0.)
R_D52130xxU24 ( 2102 2100 )  100.n
R_D52130LOADxxU24 ( 2102 0 ) COMPLEX( 390., 0.)
R_D52131xxU24 ( 2101 2100 )  100.n
R_D52131LOADxxU24 ( 2101 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU24 ( 2099 2100 )  100.n
R_D52132LOADxxU24 ( 2099 0 ) COMPLEX( 390., 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U25CCM 
R_D52101xxU25 ( 2134 2166 )  100.n
R_D52101LOADxxU25 ( 0 2166 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU25 ( 2165 2134 )  100.n
R_D52102LOADxxU25 ( 0 2165 ) COMPLEX( 390., 0.)
R_D52103xxU25 ( 2164 2134 )  100.n
R_D52103LOADxxU25 ( 0 2164 ) COMPLEX( 390., 0.)
R_D52104xxU25 ( 2163 2134 )  100.n
R_D52104LOADxxU25 ( 0 2163 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU25 ( 2162 2134 )  100.n
R_D52105LOADxxU25 ( 0 2162 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU25 ( 2161 2134 )  100.n
R_D52106LOADxxU25 ( 0 2161 ) COMPLEX( 390., 0.)
R_D52107LOADxxU25 ( 0 2159 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU25 ( 0 2160 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU25 ( 2160 2134 )  100.n
R_D52107xxU25 ( 2159 2134 )  100.n
R_D52109xxU25 ( 2158 2134 )  100.n
R_D52109LOADxxU25 ( 2158 0 ) COMPLEX( 390., 0.)
R_D52110xxU25 ( 2157 2134 )  100.n
R_D52110LOADxxU25 ( 2157 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU25 ( 2156 2134 )  100.n
R_D52111LOADxxU25 ( 2156 0 ) COMPLEX( 390., 0.)
R_D52112xxU25 ( 2155 2134 )  100.n
R_D52112LOADxxU25 ( 2155 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU25 ( 2154 2134 )  100.n
R_D52113LOADxxU25 ( 2154 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU25 ( 2153 2134 )  100.n
R_D52114LOADxxU25 ( 2153 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU25 ( 2152 2134 )  100.n
R_D52116LOADxxU25 ( 2152 0 ) COMPLEX( 390., 0.)
R_D52ExxU25 ( 548 2134 )  100.n
R_D52115xxU25 ( 2150 2134 )  100.n
R_D52115LOADxxU25 ( 2150 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU25 ( 2134 2149 )  100.n
R_D52118LOADxxU25 ( 0 2149 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU25 ( 2148 2134 )  100.n
R_D52119LOADxxU25 ( 0 2148 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU25 ( 2147 2134 )  100.n
R_D52120LOADxxU25 ( 0 2147 ) COMPLEX( 390., 0.)
R_D52121xxU25 ( 2146 2134 )  100.n
R_D52121LOADxxU25 ( 0 2146 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU25 ( 2145 2134 )  100.n
R_D52122LOADxxU25 ( 0 2145 ) COMPLEX( 390., 0.)
R_D52123xxU25 ( 2144 2134 )  100.n
R_D52123LOADxxU25 ( 0 2144 ) COMPLEX( 390., 0.)
R_D52124LOADxxU25 ( 0 2142 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU25 ( 0 2143 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU25 ( 2143 2134 )  100.n
R_D52124xxU25 ( 2142 2134 )  100.n
R_D52125xxU25 ( 2141 2134 )  100.n
R_D52125LOADxxU25 ( 2141 0 ) COMPLEX( 390., 0.)
R_D52126xxU25 ( 2140 2134 )  100.n
R_D52126LOADxxU25 ( 2140 0 ) COMPLEX( 390., 0.)
R_D52127xxU25 ( 2139 2134 )  100.n
R_D52127LOADxxU25 ( 2139 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU25 ( 2138 2134 )  100.n
R_D52128LOADxxU25 ( 2138 0 ) COMPLEX( 390., 0.)
R_D52129xxU25 ( 2137 2134 )  100.n
R_D52129LOADxxU25 ( 2137 0 ) COMPLEX( 390., 0.)
R_D52130xxU25 ( 2136 2134 )  100.n
R_D52130LOADxxU25 ( 2136 0 ) COMPLEX( 390., 0.)
R_D52131xxU25 ( 2135 2134 )  100.n
R_D52131LOADxxU25 ( 2135 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU25 ( 2133 2134 )  100.n
R_D52132LOADxxU25 ( 2133 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U26CCM 
R_D52101xxU26 ( 2168 2200 )  100.n
R_D52101LOADxxU26 ( 0 2200 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU26 ( 2199 2168 )  100.n
R_D52102LOADxxU26 ( 0 2199 ) COMPLEX( 390., 0.)
R_D52103xxU26 ( 2198 2168 )  100.n
R_D52103LOADxxU26 ( 0 2198 ) COMPLEX( 390., 0.)
R_D52104xxU26 ( 2197 2168 )  100.n
R_D52104LOADxxU26 ( 0 2197 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU26 ( 2196 2168 )  100.n
R_D52105LOADxxU26 ( 0 2196 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU26 ( 2195 2168 )  100.n
R_D52106LOADxxU26 ( 0 2195 ) COMPLEX( 390., 0.)
R_D52107LOADxxU26 ( 0 2193 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU26 ( 0 2194 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU26 ( 2194 2168 )  100.n
R_D52107xxU26 ( 2193 2168 )  100.n
R_D52109xxU26 ( 2192 2168 )  100.n
R_D52109LOADxxU26 ( 2192 0 ) COMPLEX( 390., 0.)
R_D52110xxU26 ( 2191 2168 )  100.n
R_D52110LOADxxU26 ( 2191 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU26 ( 2190 2168 )  100.n
R_D52111LOADxxU26 ( 2190 0 ) COMPLEX( 390., 0.)
R_D52112xxU26 ( 2189 2168 )  100.n
R_D52112LOADxxU26 ( 2189 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU26 ( 2188 2168 )  100.n
R_D52113LOADxxU26 ( 2188 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU26 ( 2187 2168 )  100.n
R_D52114LOADxxU26 ( 2187 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU26 ( 2186 2168 )  100.n
R_D52116LOADxxU26 ( 2186 0 ) COMPLEX( 390., 0.)
R_D52ExxU26 ( 550 2168 )  100.n
R_D52115xxU26 ( 2184 2168 )  100.n
R_D52115LOADxxU26 ( 2184 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU26 ( 2168 2183 )  100.n
R_D52118LOADxxU26 ( 0 2183 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU26 ( 2182 2168 )  100.n
R_D52119LOADxxU26 ( 0 2182 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU26 ( 2181 2168 )  100.n
R_D52120LOADxxU26 ( 0 2181 ) COMPLEX( 390., 0.)
R_D52121xxU26 ( 2180 2168 )  100.n
R_D52121LOADxxU26 ( 0 2180 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU26 ( 2179 2168 )  100.n
R_D52122LOADxxU26 ( 0 2179 ) COMPLEX( 390., 0.)
R_D52123xxU26 ( 2178 2168 )  100.n
R_D52123LOADxxU26 ( 0 2178 ) COMPLEX( 390., 0.)
R_D52124LOADxxU26 ( 0 2176 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU26 ( 0 2177 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU26 ( 2177 2168 )  100.n
R_D52124xxU26 ( 2176 2168 )  100.n
R_D52125xxU26 ( 2175 2168 )  100.n
R_D52125LOADxxU26 ( 2175 0 ) COMPLEX( 390., 0.)
R_D52126xxU26 ( 2174 2168 )  100.n
R_D52126LOADxxU26 ( 2174 0 ) COMPLEX( 390., 0.)
R_D52127xxU26 ( 2173 2168 )  100.n
R_D52127LOADxxU26 ( 2173 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU26 ( 2172 2168 )  100.n
R_D52128LOADxxU26 ( 2172 0 ) COMPLEX( 390., 0.)
R_D52129xxU26 ( 2171 2168 )  100.n
R_D52129LOADxxU26 ( 2171 0 ) COMPLEX( 390., 0.)
R_D52130xxU26 ( 2170 2168 )  100.n
R_D52130LOADxxU26 ( 2170 0 ) COMPLEX( 390., 0.)
R_D52131xxU26 ( 2169 2168 )  100.n
R_D52131LOADxxU26 ( 2169 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU26 ( 2167 2168 )  100.n
R_D52132LOADxxU26 ( 2167 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U27CCM 
R_D52101xxU27 ( 2202 2234 )  100.n
R_D52101LOADxxU27 ( 0 2234 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU27 ( 2233 2202 )  100.n
R_D52102LOADxxU27 ( 0 2233 ) COMPLEX( 390., 0.)
R_D52103xxU27 ( 2232 2202 )  100.n
R_D52103LOADxxU27 ( 0 2232 ) COMPLEX( 390., 0.)
R_D52104xxU27 ( 2231 2202 )  100.n
R_D52104LOADxxU27 ( 0 2231 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU27 ( 2230 2202 )  100.n
R_D52105LOADxxU27 ( 0 2230 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU27 ( 2229 2202 )  100.n
R_D52106LOADxxU27 ( 0 2229 ) COMPLEX( 390., 0.)
R_D52107LOADxxU27 ( 0 2227 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU27 ( 0 2228 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU27 ( 2228 2202 )  100.n
R_D52107xxU27 ( 2227 2202 )  100.n
R_D52109xxU27 ( 2226 2202 )  100.n
R_D52109LOADxxU27 ( 2226 0 ) COMPLEX( 390., 0.)
R_D52110xxU27 ( 2225 2202 )  100.n
R_D52110LOADxxU27 ( 2225 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU27 ( 2224 2202 )  100.n
R_D52111LOADxxU27 ( 2224 0 ) COMPLEX( 390., 0.)
R_D52112xxU27 ( 2223 2202 )  100.n
R_D52112LOADxxU27 ( 2223 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU27 ( 2222 2202 )  100.n
R_D52113LOADxxU27 ( 2222 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU27 ( 2221 2202 )  100.n
R_D52114LOADxxU27 ( 2221 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU27 ( 2220 2202 )  100.n
R_D52116LOADxxU27 ( 2220 0 ) COMPLEX( 390., 0.)
R_D52ExxU27 ( 553 2202 )  100.n
R_D52115xxU27 ( 2218 2202 )  100.n
R_D52115LOADxxU27 ( 2218 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU27 ( 2202 2217 )  100.n
R_D52118LOADxxU27 ( 0 2217 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU27 ( 2216 2202 )  100.n
R_D52119LOADxxU27 ( 0 2216 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU27 ( 2215 2202 )  100.n
R_D52120LOADxxU27 ( 0 2215 ) COMPLEX( 390., 0.)
R_D52121xxU27 ( 2214 2202 )  100.n
R_D52121LOADxxU27 ( 0 2214 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU27 ( 2213 2202 )  100.n
R_D52122LOADxxU27 ( 0 2213 ) COMPLEX( 390., 0.)
R_D52123xxU27 ( 2212 2202 )  100.n
R_D52123LOADxxU27 ( 0 2212 ) COMPLEX( 390., 0.)
R_D52124LOADxxU27 ( 0 2210 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU27 ( 0 2211 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU27 ( 2211 2202 )  100.n
R_D52124xxU27 ( 2210 2202 )  100.n
R_D52125xxU27 ( 2209 2202 )  100.n
R_D52125LOADxxU27 ( 2209 0 ) COMPLEX( 390., 0.)
R_D52126xxU27 ( 2208 2202 )  100.n
R_D52126LOADxxU27 ( 2208 0 ) COMPLEX( 390., 0.)
R_D52127xxU27 ( 2207 2202 )  100.n
R_D52127LOADxxU27 ( 2207 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU27 ( 2206 2202 )  100.n
R_D52128LOADxxU27 ( 2206 0 ) COMPLEX( 390., 0.)
R_D52129xxU27 ( 2205 2202 )  100.n
R_D52129LOADxxU27 ( 2205 0 ) COMPLEX( 390., 0.)
R_D52130xxU27 ( 2204 2202 )  100.n
R_D52130LOADxxU27 ( 2204 0 ) COMPLEX( 390., 0.)
R_D52131xxU27 ( 2203 2202 )  100.n
R_D52131LOADxxU27 ( 2203 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU27 ( 2201 2202 )  100.n
R_D52132LOADxxU27 ( 2201 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U28CCM 
R_D52101xxU28 ( 2236 2268 )  100.n
R_D52101LOADxxU28 ( 0 2268 ) COMPLEX( 2.8263,-1.8255)
R_D52102xxU28 ( 2267 2236 )  100.n
R_D52102LOADxxU28 ( 0 2267 ) COMPLEX( 390., 0.)
R_D52103xxU28 ( 2266 2236 )  100.n
R_D52103LOADxxU28 ( 0 2266 ) COMPLEX( 390., 0.)
R_D52104xxU28 ( 2265 2236 )  100.n
R_D52104LOADxxU28 ( 0 2265 ) COMPLEX( 26.6742,-17.9253)
R_D52105xxU28 ( 2264 2236 )  100.n
R_D52105LOADxxU28 ( 0 2264 ) COMPLEX( 26.6742,-17.9253)
R_D52106xxU28 ( 2263 2236 )  100.n
R_D52106LOADxxU28 ( 0 2263 ) COMPLEX( 390., 0.)
R_D52107LOADxxU28 ( 0 2261 ) COMPLEX( 13.9875,-8.6688)
R_D52108LOADxxU28 ( 0 2262 ) COMPLEX( 13.9875,-8.6688)
R_D52108xxU28 ( 2262 2236 )  100.n
R_D52107xxU28 ( 2261 2236 )  100.n
R_D52109xxU28 ( 2260 2236 )  100.n
R_D52109LOADxxU28 ( 2260 0 ) COMPLEX( 390., 0.)
R_D52110xxU28 ( 2259 2236 )  100.n
R_D52110LOADxxU28 ( 2259 0 ) COMPLEX( 8.1777,-4.4139)
R_D52111xxU28 ( 2258 2236 )  100.n
R_D52111LOADxxU28 ( 2258 0 ) COMPLEX( 390., 0.)
R_D52112xxU28 ( 2257 2236 )  100.n
R_D52112LOADxxU28 ( 2257 0 ) COMPLEX( 3.9963,-2.265)
R_D52113xxU28 ( 2256 2236 )  100.n
R_D52113LOADxxU28 ( 2256 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxU28 ( 2255 2236 )  100.n
R_D52114LOADxxU28 ( 2255 0 ) COMPLEX( 69.7374,-48.6771)
R_D52116xxU28 ( 2254 2236 )  100.n
R_D52116LOADxxU28 ( 2254 0 ) COMPLEX( 390., 0.)
R_D52ExxU28 ( 552 2236 )  100.n
R_D52115xxU28 ( 2252 2236 )  100.n
R_D52115LOADxxU28 ( 2252 0 ) COMPLEX( 69.7374,-48.6771)
R_D52118xxU28 ( 2236 2251 )  100.n
R_D52118LOADxxU28 ( 0 2251 ) COMPLEX( 1.363267K,-1.593835K)
R_D52119xxU28 ( 2250 2236 )  100.n
R_D52119LOADxxU28 ( 0 2250 ) COMPLEX( 1.363267K,-1.593835K)
R_D52120xxU28 ( 2249 2236 )  100.n
R_D52120LOADxxU28 ( 0 2249 ) COMPLEX( 390., 0.)
R_D52121xxU28 ( 2248 2236 )  100.n
R_D52121LOADxxU28 ( 0 2248 ) COMPLEX( 95.2656,-68.9712)
R_D52122xxU28 ( 2247 2236 )  100.n
R_D52122LOADxxU28 ( 0 2247 ) COMPLEX( 390., 0.)
R_D52123xxU28 ( 2246 2236 )  100.n
R_D52123LOADxxU28 ( 0 2246 ) COMPLEX( 390., 0.)
R_D52124LOADxxU28 ( 0 2244 ) COMPLEX( 176.6793,-141.7467)
R_D52117LOADxxU28 ( 0 2245 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU28 ( 2245 2236 )  100.n
R_D52124xxU28 ( 2244 2236 )  100.n
R_D52125xxU28 ( 2243 2236 )  100.n
R_D52125LOADxxU28 ( 2243 0 ) COMPLEX( 390., 0.)
R_D52126xxU28 ( 2242 2236 )  100.n
R_D52126LOADxxU28 ( 2242 0 ) COMPLEX( 390., 0.)
R_D52127xxU28 ( 2241 2236 )  100.n
R_D52127LOADxxU28 ( 2241 0 ) COMPLEX( 76.5744,-53.4492)
R_D52128xxU28 ( 2240 2236 )  100.n
R_D52128LOADxxU28 ( 2240 0 ) COMPLEX( 390., 0.)
R_D52129xxU28 ( 2239 2236 )  100.n
R_D52129LOADxxU28 ( 2239 0 ) COMPLEX( 390., 0.)
R_D52130xxU28 ( 2238 2236 )  100.n
R_D52130LOADxxU28 ( 2238 0 ) COMPLEX( 390., 0.)
R_D52131xxU28 ( 2237 2236 )  100.n
R_D52131LOADxxU28 ( 2237 0 ) COMPLEX( 220.8492,-177.1833)
R_D52132xxU28 ( 2235 2236 )  100.n
R_D52132LOADxxU28 ( 2235 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U29CCM 
R_D52101xxU29 ( 2270 2301 )  100.n
R_D52101LOADxxU29 ( 0 2301 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU29 ( 2300 2270 )  100.n
R_D52102LOADxxU29 ( 0 2300 ) COMPLEX( 390., 0.)
R_D52103xxU29 ( 2299 2270 )  100.n
R_D52103LOADxxU29 ( 0 2299 ) COMPLEX( 390., 0.)
R_D52104xxU29 ( 2298 2270 )  100.n
R_D52104LOADxxU29 ( 0 2298 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU29 ( 2297 2270 )  100.n
R_D52105LOADxxU29 ( 0 2297 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU29 ( 2296 2270 )  100.n
R_D52106LOADxxU29 ( 0 2296 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU29 ( 0 2294 ) COMPLEX( 390., 0.)
R_D52108LOADxxU29 ( 0 2295 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU29 ( 2295 2270 )  100.n
R_D52107xxU29 ( 2294 2270 )  100.n
R_D52109xxU29 ( 2293 2270 )  100.n
R_D52109LOADxxU29 ( 2293 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU29 ( 2292 2270 )  100.n
R_D52110LOADxxU29 ( 2292 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU29 ( 2291 2270 )  100.n
R_D52111LOADxxU29 ( 2291 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU29 ( 2290 2270 )  100.n
R_D52112LOADxxU29 ( 2290 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU29 ( 2289 2270 )  100.n
R_D52113LOADxxU29 ( 2289 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU29 ( 2288 2270 )  100.n
R_D52114LOADxxU29 ( 2288 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU29 ( 2287 2270 )  100.n
R_D52116LOADxxU29 ( 2287 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU29 ( 605 2270 )  100.n
R_D52115xxU29 ( 2285 2270 )  100.n
R_D52115LOADxxU29 ( 2285 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU29 ( 2270 2284 )  100.n
R_D52118LOADxxU29 ( 0 2284 ) COMPLEX( 390., 0.)
R_D52119xxU29 ( 2283 2270 )  100.n
R_D52119LOADxxU29 ( 0 2283 ) COMPLEX( 390., 0.)
R_D52120xxU29 ( 2282 2270 )  100.n
R_D52120LOADxxU29 ( 0 2282 ) COMPLEX( 390., 0.)
R_D52121xxU29 ( 2281 2270 )  100.n
R_D52121LOADxxU29 ( 0 2281 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU29 ( 2280 2270 )  100.n
R_D52122LOADxxU29 ( 0 2280 ) COMPLEX( 151.656,-121.671)
R_D52123xxU29 ( 2279 2270 )  100.n
R_D52123LOADxxU29 ( 0 2279 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU29 ( 0 2277 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU29 ( 0 2278 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU29 ( 2278 2270 )  100.n
R_D52124xxU29 ( 2277 2270 )  100.n
R_D52125xxU29 ( 2276 2270 )  100.n
R_D52125LOADxxU29 ( 2276 0 ) COMPLEX( 390., 0.)
R_D52126xxU29 ( 2275 2270 )  100.n
R_D52126LOADxxU29 ( 2275 0 ) COMPLEX( 390., 0.)
R_D52127xxU29 ( 2274 2270 )  100.n
R_D52127LOADxxU29 ( 2274 0 ) COMPLEX( 390., 0.)
R_D52128xxU29 ( 2273 2270 )  100.n
R_D52128LOADxxU29 ( 2273 0 ) COMPLEX( 390., 0.)
R_D52129xxU29 ( 2272 2270 )  100.n
R_D52129LOADxxU29 ( 2272 0 ) COMPLEX( 390., 0.)
R_D52130xxU29 ( 2271 2270 )  100.n
R_D52130LOADxxU29 ( 2271 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU29 ( 2269 2270 )  100.n
R_D52131LOADxxU29 ( 2269 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U30CCM 
R_D52101xxU30 ( 2303 2334 )  100.n
R_D52101LOADxxU30 ( 0 2334 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU30 ( 2333 2303 )  100.n
R_D52102LOADxxU30 ( 0 2333 ) COMPLEX( 390., 0.)
R_D52103xxU30 ( 2332 2303 )  100.n
R_D52103LOADxxU30 ( 0 2332 ) COMPLEX( 390., 0.)
R_D52104xxU30 ( 2331 2303 )  100.n
R_D52104LOADxxU30 ( 0 2331 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU30 ( 2330 2303 )  100.n
R_D52105LOADxxU30 ( 0 2330 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU30 ( 2329 2303 )  100.n
R_D52106LOADxxU30 ( 0 2329 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU30 ( 0 2327 ) COMPLEX( 390., 0.)
R_D52108LOADxxU30 ( 0 2328 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU30 ( 2328 2303 )  100.n
R_D52107xxU30 ( 2327 2303 )  100.n
R_D52109xxU30 ( 2326 2303 )  100.n
R_D52109LOADxxU30 ( 2326 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU30 ( 2325 2303 )  100.n
R_D52110LOADxxU30 ( 2325 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU30 ( 2324 2303 )  100.n
R_D52111LOADxxU30 ( 2324 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU30 ( 2323 2303 )  100.n
R_D52112LOADxxU30 ( 2323 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU30 ( 2322 2303 )  100.n
R_D52113LOADxxU30 ( 2322 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU30 ( 2321 2303 )  100.n
R_D52114LOADxxU30 ( 2321 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU30 ( 2320 2303 )  100.n
R_D52116LOADxxU30 ( 2320 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU30 ( 607 2303 )  100.n
R_D52115xxU30 ( 2318 2303 )  100.n
R_D52115LOADxxU30 ( 2318 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU30 ( 2303 2317 )  100.n
R_D52118LOADxxU30 ( 0 2317 ) COMPLEX( 390., 0.)
R_D52119xxU30 ( 2316 2303 )  100.n
R_D52119LOADxxU30 ( 0 2316 ) COMPLEX( 390., 0.)
R_D52120xxU30 ( 2315 2303 )  100.n
R_D52120LOADxxU30 ( 0 2315 ) COMPLEX( 390., 0.)
R_D52121xxU30 ( 2314 2303 )  100.n
R_D52121LOADxxU30 ( 0 2314 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU30 ( 2313 2303 )  100.n
R_D52122LOADxxU30 ( 0 2313 ) COMPLEX( 151.656,-121.671)
R_D52123xxU30 ( 2312 2303 )  100.n
R_D52123LOADxxU30 ( 0 2312 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU30 ( 0 2310 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU30 ( 0 2311 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU30 ( 2311 2303 )  100.n
R_D52124xxU30 ( 2310 2303 )  100.n
R_D52125xxU30 ( 2309 2303 )  100.n
R_D52125LOADxxU30 ( 2309 0 ) COMPLEX( 390., 0.)
R_D52126xxU30 ( 2308 2303 )  100.n
R_D52126LOADxxU30 ( 2308 0 ) COMPLEX( 390., 0.)
R_D52127xxU30 ( 2307 2303 )  100.n
R_D52127LOADxxU30 ( 2307 0 ) COMPLEX( 390., 0.)
R_D52128xxU30 ( 2306 2303 )  100.n
R_D52128LOADxxU30 ( 2306 0 ) COMPLEX( 390., 0.)
R_D52129xxU30 ( 2305 2303 )  100.n
R_D52129LOADxxU30 ( 2305 0 ) COMPLEX( 390., 0.)
R_D52130xxU30 ( 2304 2303 )  100.n
R_D52130LOADxxU30 ( 2304 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU30 ( 2302 2303 )  100.n
R_D52131LOADxxU30 ( 2302 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U31CCM 
R_D52101xxU31 ( 2336 2367 )  100.n
R_D52101LOADxxU31 ( 0 2367 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU31 ( 2366 2336 )  100.n
R_D52102LOADxxU31 ( 0 2366 ) COMPLEX( 390., 0.)
R_D52103xxU31 ( 2365 2336 )  100.n
R_D52103LOADxxU31 ( 0 2365 ) COMPLEX( 390., 0.)
R_D52104xxU31 ( 2364 2336 )  100.n
R_D52104LOADxxU31 ( 0 2364 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU31 ( 2363 2336 )  100.n
R_D52105LOADxxU31 ( 0 2363 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU31 ( 2362 2336 )  100.n
R_D52106LOADxxU31 ( 0 2362 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU31 ( 0 2360 ) COMPLEX( 390., 0.)
R_D52108LOADxxU31 ( 0 2361 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU31 ( 2361 2336 )  100.n
R_D52107xxU31 ( 2360 2336 )  100.n
R_D52109xxU31 ( 2359 2336 )  100.n
R_D52109LOADxxU31 ( 2359 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU31 ( 2358 2336 )  100.n
R_D52110LOADxxU31 ( 2358 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU31 ( 2357 2336 )  100.n
R_D52111LOADxxU31 ( 2357 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU31 ( 2356 2336 )  100.n
R_D52112LOADxxU31 ( 2356 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU31 ( 2355 2336 )  100.n
R_D52113LOADxxU31 ( 2355 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU31 ( 2354 2336 )  100.n
R_D52114LOADxxU31 ( 2354 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU31 ( 2353 2336 )  100.n
R_D52116LOADxxU31 ( 2353 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU31 ( 611 2336 )  100.n
R_D52115xxU31 ( 2351 2336 )  100.n
R_D52115LOADxxU31 ( 2351 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU31 ( 2336 2350 )  100.n
R_D52118LOADxxU31 ( 0 2350 ) COMPLEX( 390., 0.)
R_D52119xxU31 ( 2349 2336 )  100.n
R_D52119LOADxxU31 ( 0 2349 ) COMPLEX( 390., 0.)
R_D52120xxU31 ( 2348 2336 )  100.n
R_D52120LOADxxU31 ( 0 2348 ) COMPLEX( 390., 0.)
R_D52121xxU31 ( 2347 2336 )  100.n
R_D52121LOADxxU31 ( 0 2347 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU31 ( 2346 2336 )  100.n
R_D52122LOADxxU31 ( 0 2346 ) COMPLEX( 151.656,-121.671)
R_D52123xxU31 ( 2345 2336 )  100.n
R_D52123LOADxxU31 ( 0 2345 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU31 ( 0 2343 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU31 ( 0 2344 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU31 ( 2344 2336 )  100.n
R_D52124xxU31 ( 2343 2336 )  100.n
R_D52125xxU31 ( 2342 2336 )  100.n
R_D52125LOADxxU31 ( 2342 0 ) COMPLEX( 390., 0.)
R_D52126xxU31 ( 2341 2336 )  100.n
R_D52126LOADxxU31 ( 2341 0 ) COMPLEX( 390., 0.)
R_D52127xxU31 ( 2340 2336 )  100.n
R_D52127LOADxxU31 ( 2340 0 ) COMPLEX( 390., 0.)
R_D52128xxU31 ( 2339 2336 )  100.n
R_D52128LOADxxU31 ( 2339 0 ) COMPLEX( 390., 0.)
R_D52129xxU31 ( 2338 2336 )  100.n
R_D52129LOADxxU31 ( 2338 0 ) COMPLEX( 390., 0.)
R_D52130xxU31 ( 2337 2336 )  100.n
R_D52130LOADxxU31 ( 2337 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU31 ( 2335 2336 )  100.n
R_D52131LOADxxU31 ( 2335 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U32CCM 
R_D52101xxU32 ( 2369 2400 )  100.n
R_D52101LOADxxU32 ( 0 2400 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU32 ( 2399 2369 )  100.n
R_D52102LOADxxU32 ( 0 2399 ) COMPLEX( 390., 0.)
R_D52103xxU32 ( 2398 2369 )  100.n
R_D52103LOADxxU32 ( 0 2398 ) COMPLEX( 390., 0.)
R_D52104xxU32 ( 2397 2369 )  100.n
R_D52104LOADxxU32 ( 0 2397 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU32 ( 2396 2369 )  100.n
R_D52105LOADxxU32 ( 0 2396 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU32 ( 2395 2369 )  100.n
R_D52106LOADxxU32 ( 0 2395 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU32 ( 0 2393 ) COMPLEX( 390., 0.)
R_D52108LOADxxU32 ( 0 2394 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU32 ( 2394 2369 )  100.n
R_D52107xxU32 ( 2393 2369 )  100.n
R_D52109xxU32 ( 2392 2369 )  100.n
R_D52109LOADxxU32 ( 2392 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU32 ( 2391 2369 )  100.n
R_D52110LOADxxU32 ( 2391 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU32 ( 2390 2369 )  100.n
R_D52111LOADxxU32 ( 2390 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU32 ( 2389 2369 )  100.n
R_D52112LOADxxU32 ( 2389 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU32 ( 2388 2369 )  100.n
R_D52113LOADxxU32 ( 2388 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU32 ( 2387 2369 )  100.n
R_D52114LOADxxU32 ( 2387 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU32 ( 2386 2369 )  100.n
R_D52116LOADxxU32 ( 2386 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU32 ( 610 2369 )  100.n
R_D52115xxU32 ( 2384 2369 )  100.n
R_D52115LOADxxU32 ( 2384 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU32 ( 2369 2383 )  100.n
R_D52118LOADxxU32 ( 0 2383 ) COMPLEX( 390., 0.)
R_D52119xxU32 ( 2382 2369 )  100.n
R_D52119LOADxxU32 ( 0 2382 ) COMPLEX( 390., 0.)
R_D52120xxU32 ( 2381 2369 )  100.n
R_D52120LOADxxU32 ( 0 2381 ) COMPLEX( 390., 0.)
R_D52121xxU32 ( 2380 2369 )  100.n
R_D52121LOADxxU32 ( 0 2380 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU32 ( 2379 2369 )  100.n
R_D52122LOADxxU32 ( 0 2379 ) COMPLEX( 151.656,-121.671)
R_D52123xxU32 ( 2378 2369 )  100.n
R_D52123LOADxxU32 ( 0 2378 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU32 ( 0 2376 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU32 ( 0 2377 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU32 ( 2377 2369 )  100.n
R_D52124xxU32 ( 2376 2369 )  100.n
R_D52125xxU32 ( 2375 2369 )  100.n
R_D52125LOADxxU32 ( 2375 0 ) COMPLEX( 390., 0.)
R_D52126xxU32 ( 2374 2369 )  100.n
R_D52126LOADxxU32 ( 2374 0 ) COMPLEX( 390., 0.)
R_D52127xxU32 ( 2373 2369 )  100.n
R_D52127LOADxxU32 ( 2373 0 ) COMPLEX( 390., 0.)
R_D52128xxU32 ( 2372 2369 )  100.n
R_D52128LOADxxU32 ( 2372 0 ) COMPLEX( 390., 0.)
R_D52129xxU32 ( 2371 2369 )  100.n
R_D52129LOADxxU32 ( 2371 0 ) COMPLEX( 390., 0.)
R_D52130xxU32 ( 2370 2369 )  100.n
R_D52130LOADxxU32 ( 2370 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU32 ( 2368 2369 )  100.n
R_D52131LOADxxU32 ( 2368 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U33CCM 
R_D52101xxU33 ( 2402 2433 )  100.n
R_D52101LOADxxU33 ( 0 2433 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU33 ( 2432 2402 )  100.n
R_D52102LOADxxU33 ( 0 2432 ) COMPLEX( 390., 0.)
R_D52103xxU33 ( 2431 2402 )  100.n
R_D52103LOADxxU33 ( 0 2431 ) COMPLEX( 390., 0.)
R_D52104xxU33 ( 2430 2402 )  100.n
R_D52104LOADxxU33 ( 0 2430 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU33 ( 2429 2402 )  100.n
R_D52105LOADxxU33 ( 0 2429 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU33 ( 2428 2402 )  100.n
R_D52106LOADxxU33 ( 0 2428 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU33 ( 0 2426 ) COMPLEX( 390., 0.)
R_D52108LOADxxU33 ( 0 2427 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU33 ( 2427 2402 )  100.n
R_D52107xxU33 ( 2426 2402 )  100.n
R_D52109xxU33 ( 2425 2402 )  100.n
R_D52109LOADxxU33 ( 2425 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU33 ( 2424 2402 )  100.n
R_D52110LOADxxU33 ( 2424 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU33 ( 2423 2402 )  100.n
R_D52111LOADxxU33 ( 2423 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU33 ( 2422 2402 )  100.n
R_D52112LOADxxU33 ( 2422 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU33 ( 2421 2402 )  100.n
R_D52113LOADxxU33 ( 2421 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU33 ( 2420 2402 )  100.n
R_D52114LOADxxU33 ( 2420 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU33 ( 2419 2402 )  100.n
R_D52116LOADxxU33 ( 2419 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU33 ( 489 2402 )  100.n
R_D52115xxU33 ( 2417 2402 )  100.n
R_D52115LOADxxU33 ( 2417 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU33 ( 2402 2416 )  100.n
R_D52118LOADxxU33 ( 0 2416 ) COMPLEX( 390., 0.)
R_D52119xxU33 ( 2415 2402 )  100.n
R_D52119LOADxxU33 ( 0 2415 ) COMPLEX( 390., 0.)
R_D52120xxU33 ( 2414 2402 )  100.n
R_D52120LOADxxU33 ( 0 2414 ) COMPLEX( 390., 0.)
R_D52121xxU33 ( 2413 2402 )  100.n
R_D52121LOADxxU33 ( 0 2413 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU33 ( 2412 2402 )  100.n
R_D52122LOADxxU33 ( 0 2412 ) COMPLEX( 151.656,-121.671)
R_D52123xxU33 ( 2411 2402 )  100.n
R_D52123LOADxxU33 ( 0 2411 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU33 ( 0 2409 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU33 ( 0 2410 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU33 ( 2410 2402 )  100.n
R_D52124xxU33 ( 2409 2402 )  100.n
R_D52125xxU33 ( 2408 2402 )  100.n
R_D52125LOADxxU33 ( 2408 0 ) COMPLEX( 390., 0.)
R_D52126xxU33 ( 2407 2402 )  100.n
R_D52126LOADxxU33 ( 2407 0 ) COMPLEX( 390., 0.)
R_D52127xxU33 ( 2406 2402 )  100.n
R_D52127LOADxxU33 ( 2406 0 ) COMPLEX( 390., 0.)
R_D52128xxU33 ( 2405 2402 )  100.n
R_D52128LOADxxU33 ( 2405 0 ) COMPLEX( 390., 0.)
R_D52129xxU33 ( 2404 2402 )  100.n
R_D52129LOADxxU33 ( 2404 0 ) COMPLEX( 390., 0.)
R_D52130xxU33 ( 2403 2402 )  100.n
R_D52130LOADxxU33 ( 2403 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU33 ( 2401 2402 )  100.n
R_D52131LOADxxU33 ( 2401 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U34CCM 
R_D52101xxU34 ( 2435 2466 )  100.n
R_D52101LOADxxU34 ( 0 2466 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU34 ( 2465 2435 )  100.n
R_D52102LOADxxU34 ( 0 2465 ) COMPLEX( 390., 0.)
R_D52103xxU34 ( 2464 2435 )  100.n
R_D52103LOADxxU34 ( 0 2464 ) COMPLEX( 390., 0.)
R_D52104xxU34 ( 2463 2435 )  100.n
R_D52104LOADxxU34 ( 0 2463 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU34 ( 2462 2435 )  100.n
R_D52105LOADxxU34 ( 0 2462 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU34 ( 2461 2435 )  100.n
R_D52106LOADxxU34 ( 0 2461 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU34 ( 0 2459 ) COMPLEX( 390., 0.)
R_D52108LOADxxU34 ( 0 2460 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU34 ( 2460 2435 )  100.n
R_D52107xxU34 ( 2459 2435 )  100.n
R_D52109xxU34 ( 2458 2435 )  100.n
R_D52109LOADxxU34 ( 2458 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU34 ( 2457 2435 )  100.n
R_D52110LOADxxU34 ( 2457 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU34 ( 2456 2435 )  100.n
R_D52111LOADxxU34 ( 2456 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU34 ( 2455 2435 )  100.n
R_D52112LOADxxU34 ( 2455 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU34 ( 2454 2435 )  100.n
R_D52113LOADxxU34 ( 2454 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU34 ( 2453 2435 )  100.n
R_D52114LOADxxU34 ( 2453 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU34 ( 2452 2435 )  100.n
R_D52116LOADxxU34 ( 2452 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU34 ( 491 2435 )  100.n
R_D52115xxU34 ( 2450 2435 )  100.n
R_D52115LOADxxU34 ( 2450 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU34 ( 2435 2449 )  100.n
R_D52118LOADxxU34 ( 0 2449 ) COMPLEX( 390., 0.)
R_D52119xxU34 ( 2448 2435 )  100.n
R_D52119LOADxxU34 ( 0 2448 ) COMPLEX( 390., 0.)
R_D52120xxU34 ( 2447 2435 )  100.n
R_D52120LOADxxU34 ( 0 2447 ) COMPLEX( 390., 0.)
R_D52121xxU34 ( 2446 2435 )  100.n
R_D52121LOADxxU34 ( 0 2446 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU34 ( 2445 2435 )  100.n
R_D52122LOADxxU34 ( 0 2445 ) COMPLEX( 151.656,-121.671)
R_D52123xxU34 ( 2444 2435 )  100.n
R_D52123LOADxxU34 ( 0 2444 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU34 ( 0 2442 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU34 ( 0 2443 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU34 ( 2443 2435 )  100.n
R_D52124xxU34 ( 2442 2435 )  100.n
R_D52125xxU34 ( 2441 2435 )  100.n
R_D52125LOADxxU34 ( 2441 0 ) COMPLEX( 390., 0.)
R_D52126xxU34 ( 2440 2435 )  100.n
R_D52126LOADxxU34 ( 2440 0 ) COMPLEX( 390., 0.)
R_D52127xxU34 ( 2439 2435 )  100.n
R_D52127LOADxxU34 ( 2439 0 ) COMPLEX( 390., 0.)
R_D52128xxU34 ( 2438 2435 )  100.n
R_D52128LOADxxU34 ( 2438 0 ) COMPLEX( 390., 0.)
R_D52129xxU34 ( 2437 2435 )  100.n
R_D52129LOADxxU34 ( 2437 0 ) COMPLEX( 390., 0.)
R_D52130xxU34 ( 2436 2435 )  100.n
R_D52130LOADxxU34 ( 2436 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU34 ( 2434 2435 )  100.n
R_D52131LOADxxU34 ( 2434 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U35CCM 
R_D52101xxU35 ( 2468 2499 )  100.n
R_D52101LOADxxU35 ( 0 2499 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU35 ( 2498 2468 )  100.n
R_D52102LOADxxU35 ( 0 2498 ) COMPLEX( 390., 0.)
R_D52103xxU35 ( 2497 2468 )  100.n
R_D52103LOADxxU35 ( 0 2497 ) COMPLEX( 390., 0.)
R_D52104xxU35 ( 2496 2468 )  100.n
R_D52104LOADxxU35 ( 0 2496 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU35 ( 2495 2468 )  100.n
R_D52105LOADxxU35 ( 0 2495 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU35 ( 2494 2468 )  100.n
R_D52106LOADxxU35 ( 0 2494 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU35 ( 0 2492 ) COMPLEX( 390., 0.)
R_D52108LOADxxU35 ( 0 2493 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU35 ( 2493 2468 )  100.n
R_D52107xxU35 ( 2492 2468 )  100.n
R_D52109xxU35 ( 2491 2468 )  100.n
R_D52109LOADxxU35 ( 2491 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU35 ( 2490 2468 )  100.n
R_D52110LOADxxU35 ( 2490 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU35 ( 2489 2468 )  100.n
R_D52111LOADxxU35 ( 2489 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU35 ( 2488 2468 )  100.n
R_D52112LOADxxU35 ( 2488 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU35 ( 2487 2468 )  100.n
R_D52113LOADxxU35 ( 2487 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU35 ( 2486 2468 )  100.n
R_D52114LOADxxU35 ( 2486 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU35 ( 2485 2468 )  100.n
R_D52116LOADxxU35 ( 2485 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU35 ( 495 2468 )  100.n
R_D52115xxU35 ( 2483 2468 )  100.n
R_D52115LOADxxU35 ( 2483 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU35 ( 2468 2482 )  100.n
R_D52118LOADxxU35 ( 0 2482 ) COMPLEX( 390., 0.)
R_D52119xxU35 ( 2481 2468 )  100.n
R_D52119LOADxxU35 ( 0 2481 ) COMPLEX( 390., 0.)
R_D52120xxU35 ( 2480 2468 )  100.n
R_D52120LOADxxU35 ( 0 2480 ) COMPLEX( 390., 0.)
R_D52121xxU35 ( 2479 2468 )  100.n
R_D52121LOADxxU35 ( 0 2479 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU35 ( 2478 2468 )  100.n
R_D52122LOADxxU35 ( 0 2478 ) COMPLEX( 151.656,-121.671)
R_D52123xxU35 ( 2477 2468 )  100.n
R_D52123LOADxxU35 ( 0 2477 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU35 ( 0 2475 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU35 ( 0 2476 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU35 ( 2476 2468 )  100.n
R_D52124xxU35 ( 2475 2468 )  100.n
R_D52125xxU35 ( 2474 2468 )  100.n
R_D52125LOADxxU35 ( 2474 0 ) COMPLEX( 390., 0.)
R_D52126xxU35 ( 2473 2468 )  100.n
R_D52126LOADxxU35 ( 2473 0 ) COMPLEX( 390., 0.)
R_D52127xxU35 ( 2472 2468 )  100.n
R_D52127LOADxxU35 ( 2472 0 ) COMPLEX( 390., 0.)
R_D52128xxU35 ( 2471 2468 )  100.n
R_D52128LOADxxU35 ( 2471 0 ) COMPLEX( 390., 0.)
R_D52129xxU35 ( 2470 2468 )  100.n
R_D52129LOADxxU35 ( 2470 0 ) COMPLEX( 390., 0.)
R_D52130xxU35 ( 2469 2468 )  100.n
R_D52130LOADxxU35 ( 2469 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU35 ( 2467 2468 )  100.n
R_D52131LOADxxU35 ( 2467 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U36CCM 
R_D52101xxU36 ( 2501 2532 )  100.n
R_D52101LOADxxU36 ( 0 2532 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU36 ( 2531 2501 )  100.n
R_D52102LOADxxU36 ( 0 2531 ) COMPLEX( 390., 0.)
R_D52103xxU36 ( 2530 2501 )  100.n
R_D52103LOADxxU36 ( 0 2530 ) COMPLEX( 390., 0.)
R_D52104xxU36 ( 2529 2501 )  100.n
R_D52104LOADxxU36 ( 0 2529 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU36 ( 2528 2501 )  100.n
R_D52105LOADxxU36 ( 0 2528 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU36 ( 2527 2501 )  100.n
R_D52106LOADxxU36 ( 0 2527 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU36 ( 0 2525 ) COMPLEX( 390., 0.)
R_D52108LOADxxU36 ( 0 2526 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU36 ( 2526 2501 )  100.n
R_D52107xxU36 ( 2525 2501 )  100.n
R_D52109xxU36 ( 2524 2501 )  100.n
R_D52109LOADxxU36 ( 2524 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU36 ( 2523 2501 )  100.n
R_D52110LOADxxU36 ( 2523 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU36 ( 2522 2501 )  100.n
R_D52111LOADxxU36 ( 2522 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU36 ( 2521 2501 )  100.n
R_D52112LOADxxU36 ( 2521 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU36 ( 2520 2501 )  100.n
R_D52113LOADxxU36 ( 2520 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU36 ( 2519 2501 )  100.n
R_D52114LOADxxU36 ( 2519 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU36 ( 2518 2501 )  100.n
R_D52116LOADxxU36 ( 2518 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU36 ( 494 2501 )  100.n
R_D52115xxU36 ( 2516 2501 )  100.n
R_D52115LOADxxU36 ( 2516 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU36 ( 2501 2515 )  100.n
R_D52118LOADxxU36 ( 0 2515 ) COMPLEX( 390., 0.)
R_D52119xxU36 ( 2514 2501 )  100.n
R_D52119LOADxxU36 ( 0 2514 ) COMPLEX( 390., 0.)
R_D52120xxU36 ( 2513 2501 )  100.n
R_D52120LOADxxU36 ( 0 2513 ) COMPLEX( 390., 0.)
R_D52121xxU36 ( 2512 2501 )  100.n
R_D52121LOADxxU36 ( 0 2512 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU36 ( 2511 2501 )  100.n
R_D52122LOADxxU36 ( 0 2511 ) COMPLEX( 151.656,-121.671)
R_D52123xxU36 ( 2510 2501 )  100.n
R_D52123LOADxxU36 ( 0 2510 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU36 ( 0 2508 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU36 ( 0 2509 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU36 ( 2509 2501 )  100.n
R_D52124xxU36 ( 2508 2501 )  100.n
R_D52125xxU36 ( 2507 2501 )  100.n
R_D52125LOADxxU36 ( 2507 0 ) COMPLEX( 390., 0.)
R_D52126xxU36 ( 2506 2501 )  100.n
R_D52126LOADxxU36 ( 2506 0 ) COMPLEX( 390., 0.)
R_D52127xxU36 ( 2505 2501 )  100.n
R_D52127LOADxxU36 ( 2505 0 ) COMPLEX( 390., 0.)
R_D52128xxU36 ( 2504 2501 )  100.n
R_D52128LOADxxU36 ( 2504 0 ) COMPLEX( 390., 0.)
R_D52129xxU36 ( 2503 2501 )  100.n
R_D52129LOADxxU36 ( 2503 0 ) COMPLEX( 390., 0.)
R_D52130xxU36 ( 2502 2501 )  100.n
R_D52130LOADxxU36 ( 2502 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU36 ( 2500 2501 )  100.n
R_D52131LOADxxU36 ( 2500 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U37CCM 
R_D52101xxU37 ( 2534 2565 )  100.n
R_D52101LOADxxU37 ( 0 2565 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU37 ( 2564 2534 )  100.n
R_D52102LOADxxU37 ( 0 2564 ) COMPLEX( 390., 0.)
R_D52103xxU37 ( 2563 2534 )  100.n
R_D52103LOADxxU37 ( 0 2563 ) COMPLEX( 390., 0.)
R_D52104xxU37 ( 2562 2534 )  100.n
R_D52104LOADxxU37 ( 0 2562 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU37 ( 2561 2534 )  100.n
R_D52105LOADxxU37 ( 0 2561 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU37 ( 2560 2534 )  100.n
R_D52106LOADxxU37 ( 0 2560 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU37 ( 0 2558 ) COMPLEX( 390., 0.)
R_D52108LOADxxU37 ( 0 2559 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU37 ( 2559 2534 )  100.n
R_D52107xxU37 ( 2558 2534 )  100.n
R_D52109xxU37 ( 2557 2534 )  100.n
R_D52109LOADxxU37 ( 2557 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU37 ( 2556 2534 )  100.n
R_D52110LOADxxU37 ( 2556 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU37 ( 2555 2534 )  100.n
R_D52111LOADxxU37 ( 2555 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU37 ( 2554 2534 )  100.n
R_D52112LOADxxU37 ( 2554 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU37 ( 2553 2534 )  100.n
R_D52113LOADxxU37 ( 2553 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU37 ( 2552 2534 )  100.n
R_D52114LOADxxU37 ( 2552 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU37 ( 2551 2534 )  100.n
R_D52116LOADxxU37 ( 2551 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU37 ( 478 2534 )  100.n
R_D52115xxU37 ( 2549 2534 )  100.n
R_D52115LOADxxU37 ( 2549 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU37 ( 2534 2548 )  100.n
R_D52118LOADxxU37 ( 0 2548 ) COMPLEX( 390., 0.)
R_D52119xxU37 ( 2547 2534 )  100.n
R_D52119LOADxxU37 ( 0 2547 ) COMPLEX( 390., 0.)
R_D52120xxU37 ( 2546 2534 )  100.n
R_D52120LOADxxU37 ( 0 2546 ) COMPLEX( 390., 0.)
R_D52121xxU37 ( 2545 2534 )  100.n
R_D52121LOADxxU37 ( 0 2545 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU37 ( 2544 2534 )  100.n
R_D52122LOADxxU37 ( 0 2544 ) COMPLEX( 151.656,-121.671)
R_D52123xxU37 ( 2543 2534 )  100.n
R_D52123LOADxxU37 ( 0 2543 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU37 ( 0 2541 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU37 ( 0 2542 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU37 ( 2542 2534 )  100.n
R_D52124xxU37 ( 2541 2534 )  100.n
R_D52125xxU37 ( 2540 2534 )  100.n
R_D52125LOADxxU37 ( 2540 0 ) COMPLEX( 390., 0.)
R_D52126xxU37 ( 2539 2534 )  100.n
R_D52126LOADxxU37 ( 2539 0 ) COMPLEX( 390., 0.)
R_D52127xxU37 ( 2538 2534 )  100.n
R_D52127LOADxxU37 ( 2538 0 ) COMPLEX( 390., 0.)
R_D52128xxU37 ( 2537 2534 )  100.n
R_D52128LOADxxU37 ( 2537 0 ) COMPLEX( 390., 0.)
R_D52129xxU37 ( 2536 2534 )  100.n
R_D52129LOADxxU37 ( 2536 0 ) COMPLEX( 390., 0.)
R_D52130xxU37 ( 2535 2534 )  100.n
R_D52130LOADxxU37 ( 2535 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU37 ( 2533 2534 )  100.n
R_D52131LOADxxU37 ( 2533 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U38CCM 
R_D52101xxU38 ( 2567 2598 )  100.n
R_D52101LOADxxU38 ( 0 2598 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU38 ( 2597 2567 )  100.n
R_D52102LOADxxU38 ( 0 2597 ) COMPLEX( 390., 0.)
R_D52103xxU38 ( 2596 2567 )  100.n
R_D52103LOADxxU38 ( 0 2596 ) COMPLEX( 390., 0.)
R_D52104xxU38 ( 2595 2567 )  100.n
R_D52104LOADxxU38 ( 0 2595 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU38 ( 2594 2567 )  100.n
R_D52105LOADxxU38 ( 0 2594 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU38 ( 2593 2567 )  100.n
R_D52106LOADxxU38 ( 0 2593 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU38 ( 0 2591 ) COMPLEX( 390., 0.)
R_D52108LOADxxU38 ( 0 2592 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU38 ( 2592 2567 )  100.n
R_D52107xxU38 ( 2591 2567 )  100.n
R_D52109xxU38 ( 2590 2567 )  100.n
R_D52109LOADxxU38 ( 2590 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU38 ( 2589 2567 )  100.n
R_D52110LOADxxU38 ( 2589 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU38 ( 2588 2567 )  100.n
R_D52111LOADxxU38 ( 2588 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU38 ( 2587 2567 )  100.n
R_D52112LOADxxU38 ( 2587 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU38 ( 2586 2567 )  100.n
R_D52113LOADxxU38 ( 2586 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU38 ( 2585 2567 )  100.n
R_D52114LOADxxU38 ( 2585 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU38 ( 2584 2567 )  100.n
R_D52116LOADxxU38 ( 2584 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU38 ( 480 2567 )  100.n
R_D52115xxU38 ( 2582 2567 )  100.n
R_D52115LOADxxU38 ( 2582 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU38 ( 2567 2581 )  100.n
R_D52118LOADxxU38 ( 0 2581 ) COMPLEX( 390., 0.)
R_D52119xxU38 ( 2580 2567 )  100.n
R_D52119LOADxxU38 ( 0 2580 ) COMPLEX( 390., 0.)
R_D52120xxU38 ( 2579 2567 )  100.n
R_D52120LOADxxU38 ( 0 2579 ) COMPLEX( 390., 0.)
R_D52121xxU38 ( 2578 2567 )  100.n
R_D52121LOADxxU38 ( 0 2578 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU38 ( 2577 2567 )  100.n
R_D52122LOADxxU38 ( 0 2577 ) COMPLEX( 151.656,-121.671)
R_D52123xxU38 ( 2576 2567 )  100.n
R_D52123LOADxxU38 ( 0 2576 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU38 ( 0 2574 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU38 ( 0 2575 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU38 ( 2575 2567 )  100.n
R_D52124xxU38 ( 2574 2567 )  100.n
R_D52125xxU38 ( 2573 2567 )  100.n
R_D52125LOADxxU38 ( 2573 0 ) COMPLEX( 390., 0.)
R_D52126xxU38 ( 2572 2567 )  100.n
R_D52126LOADxxU38 ( 2572 0 ) COMPLEX( 390., 0.)
R_D52127xxU38 ( 2571 2567 )  100.n
R_D52127LOADxxU38 ( 2571 0 ) COMPLEX( 390., 0.)
R_D52128xxU38 ( 2570 2567 )  100.n
R_D52128LOADxxU38 ( 2570 0 ) COMPLEX( 390., 0.)
R_D52129xxU38 ( 2569 2567 )  100.n
R_D52129LOADxxU38 ( 2569 0 ) COMPLEX( 390., 0.)
R_D52130xxU38 ( 2568 2567 )  100.n
R_D52130LOADxxU38 ( 2568 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU38 ( 2566 2567 )  100.n
R_D52131LOADxxU38 ( 2566 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U39CCM 
R_D52101xxU39 ( 2600 2631 )  100.n
R_D52101LOADxxU39 ( 0 2631 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU39 ( 2630 2600 )  100.n
R_D52102LOADxxU39 ( 0 2630 ) COMPLEX( 390., 0.)
R_D52103xxU39 ( 2629 2600 )  100.n
R_D52103LOADxxU39 ( 0 2629 ) COMPLEX( 390., 0.)
R_D52104xxU39 ( 2628 2600 )  100.n
R_D52104LOADxxU39 ( 0 2628 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU39 ( 2627 2600 )  100.n
R_D52105LOADxxU39 ( 0 2627 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU39 ( 2626 2600 )  100.n
R_D52106LOADxxU39 ( 0 2626 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU39 ( 0 2624 ) COMPLEX( 390., 0.)
R_D52108LOADxxU39 ( 0 2625 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU39 ( 2625 2600 )  100.n
R_D52107xxU39 ( 2624 2600 )  100.n
R_D52109xxU39 ( 2623 2600 )  100.n
R_D52109LOADxxU39 ( 2623 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU39 ( 2622 2600 )  100.n
R_D52110LOADxxU39 ( 2622 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU39 ( 2621 2600 )  100.n
R_D52111LOADxxU39 ( 2621 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU39 ( 2620 2600 )  100.n
R_D52112LOADxxU39 ( 2620 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU39 ( 2619 2600 )  100.n
R_D52113LOADxxU39 ( 2619 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU39 ( 2618 2600 )  100.n
R_D52114LOADxxU39 ( 2618 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU39 ( 2617 2600 )  100.n
R_D52116LOADxxU39 ( 2617 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU39 ( 484 2600 )  100.n
R_D52115xxU39 ( 2615 2600 )  100.n
R_D52115LOADxxU39 ( 2615 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU39 ( 2600 2614 )  100.n
R_D52118LOADxxU39 ( 0 2614 ) COMPLEX( 390., 0.)
R_D52119xxU39 ( 2613 2600 )  100.n
R_D52119LOADxxU39 ( 0 2613 ) COMPLEX( 390., 0.)
R_D52120xxU39 ( 2612 2600 )  100.n
R_D52120LOADxxU39 ( 0 2612 ) COMPLEX( 390., 0.)
R_D52121xxU39 ( 2611 2600 )  100.n
R_D52121LOADxxU39 ( 0 2611 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU39 ( 2610 2600 )  100.n
R_D52122LOADxxU39 ( 0 2610 ) COMPLEX( 151.656,-121.671)
R_D52123xxU39 ( 2609 2600 )  100.n
R_D52123LOADxxU39 ( 0 2609 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU39 ( 0 2607 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU39 ( 0 2608 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU39 ( 2608 2600 )  100.n
R_D52124xxU39 ( 2607 2600 )  100.n
R_D52125xxU39 ( 2606 2600 )  100.n
R_D52125LOADxxU39 ( 2606 0 ) COMPLEX( 390., 0.)
R_D52126xxU39 ( 2605 2600 )  100.n
R_D52126LOADxxU39 ( 2605 0 ) COMPLEX( 390., 0.)
R_D52127xxU39 ( 2604 2600 )  100.n
R_D52127LOADxxU39 ( 2604 0 ) COMPLEX( 390., 0.)
R_D52128xxU39 ( 2603 2600 )  100.n
R_D52128LOADxxU39 ( 2603 0 ) COMPLEX( 390., 0.)
R_D52129xxU39 ( 2602 2600 )  100.n
R_D52129LOADxxU39 ( 2602 0 ) COMPLEX( 390., 0.)
R_D52130xxU39 ( 2601 2600 )  100.n
R_D52130LOADxxU39 ( 2601 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU39 ( 2599 2600 )  100.n
R_D52131LOADxxU39 ( 2599 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U40CCM 
R_D52101xxU40 ( 2633 2664 )  100.n
R_D52101LOADxxU40 ( 0 2664 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU40 ( 2663 2633 )  100.n
R_D52102LOADxxU40 ( 0 2663 ) COMPLEX( 390., 0.)
R_D52103xxU40 ( 2662 2633 )  100.n
R_D52103LOADxxU40 ( 0 2662 ) COMPLEX( 390., 0.)
R_D52104xxU40 ( 2661 2633 )  100.n
R_D52104LOADxxU40 ( 0 2661 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU40 ( 2660 2633 )  100.n
R_D52105LOADxxU40 ( 0 2660 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU40 ( 2659 2633 )  100.n
R_D52106LOADxxU40 ( 0 2659 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU40 ( 0 2657 ) COMPLEX( 390., 0.)
R_D52108LOADxxU40 ( 0 2658 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU40 ( 2658 2633 )  100.n
R_D52107xxU40 ( 2657 2633 )  100.n
R_D52109xxU40 ( 2656 2633 )  100.n
R_D52109LOADxxU40 ( 2656 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU40 ( 2655 2633 )  100.n
R_D52110LOADxxU40 ( 2655 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU40 ( 2654 2633 )  100.n
R_D52111LOADxxU40 ( 2654 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU40 ( 2653 2633 )  100.n
R_D52112LOADxxU40 ( 2653 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU40 ( 2652 2633 )  100.n
R_D52113LOADxxU40 ( 2652 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU40 ( 2651 2633 )  100.n
R_D52114LOADxxU40 ( 2651 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU40 ( 2650 2633 )  100.n
R_D52116LOADxxU40 ( 2650 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU40 ( 483 2633 )  100.n
R_D52115xxU40 ( 2648 2633 )  100.n
R_D52115LOADxxU40 ( 2648 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU40 ( 2633 2647 )  100.n
R_D52118LOADxxU40 ( 0 2647 ) COMPLEX( 390., 0.)
R_D52119xxU40 ( 2646 2633 )  100.n
R_D52119LOADxxU40 ( 0 2646 ) COMPLEX( 390., 0.)
R_D52120xxU40 ( 2645 2633 )  100.n
R_D52120LOADxxU40 ( 0 2645 ) COMPLEX( 390., 0.)
R_D52121xxU40 ( 2644 2633 )  100.n
R_D52121LOADxxU40 ( 0 2644 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU40 ( 2643 2633 )  100.n
R_D52122LOADxxU40 ( 0 2643 ) COMPLEX( 151.656,-121.671)
R_D52123xxU40 ( 2642 2633 )  100.n
R_D52123LOADxxU40 ( 0 2642 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU40 ( 0 2640 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU40 ( 0 2641 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU40 ( 2641 2633 )  100.n
R_D52124xxU40 ( 2640 2633 )  100.n
R_D52125xxU40 ( 2639 2633 )  100.n
R_D52125LOADxxU40 ( 2639 0 ) COMPLEX( 390., 0.)
R_D52126xxU40 ( 2638 2633 )  100.n
R_D52126LOADxxU40 ( 2638 0 ) COMPLEX( 390., 0.)
R_D52127xxU40 ( 2637 2633 )  100.n
R_D52127LOADxxU40 ( 2637 0 ) COMPLEX( 390., 0.)
R_D52128xxU40 ( 2636 2633 )  100.n
R_D52128LOADxxU40 ( 2636 0 ) COMPLEX( 390., 0.)
R_D52129xxU40 ( 2635 2633 )  100.n
R_D52129LOADxxU40 ( 2635 0 ) COMPLEX( 390., 0.)
R_D52130xxU40 ( 2634 2633 )  100.n
R_D52130LOADxxU40 ( 2634 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU40 ( 2632 2633 )  100.n
R_D52131LOADxxU40 ( 2632 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U41CCM 
R_D52101xxU41 ( 2666 2697 )  100.n
R_D52101LOADxxU41 ( 0 2697 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU41 ( 2696 2666 )  100.n
R_D52102LOADxxU41 ( 0 2696 ) COMPLEX( 390., 0.)
R_D52103xxU41 ( 2695 2666 )  100.n
R_D52103LOADxxU41 ( 0 2695 ) COMPLEX( 390., 0.)
R_D52104xxU41 ( 2694 2666 )  100.n
R_D52104LOADxxU41 ( 0 2694 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU41 ( 2693 2666 )  100.n
R_D52105LOADxxU41 ( 0 2693 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU41 ( 2692 2666 )  100.n
R_D52106LOADxxU41 ( 0 2692 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU41 ( 0 2690 ) COMPLEX( 390., 0.)
R_D52108LOADxxU41 ( 0 2691 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU41 ( 2691 2666 )  100.n
R_D52107xxU41 ( 2690 2666 )  100.n
R_D52109xxU41 ( 2689 2666 )  100.n
R_D52109LOADxxU41 ( 2689 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU41 ( 2688 2666 )  100.n
R_D52110LOADxxU41 ( 2688 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU41 ( 2687 2666 )  100.n
R_D52111LOADxxU41 ( 2687 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU41 ( 2686 2666 )  100.n
R_D52112LOADxxU41 ( 2686 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU41 ( 2685 2666 )  100.n
R_D52113LOADxxU41 ( 2685 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU41 ( 2684 2666 )  100.n
R_D52114LOADxxU41 ( 2684 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU41 ( 2683 2666 )  100.n
R_D52116LOADxxU41 ( 2683 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU41 ( 536 2666 )  100.n
R_D52115xxU41 ( 2681 2666 )  100.n
R_D52115LOADxxU41 ( 2681 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU41 ( 2666 2680 )  100.n
R_D52118LOADxxU41 ( 0 2680 ) COMPLEX( 390., 0.)
R_D52119xxU41 ( 2679 2666 )  100.n
R_D52119LOADxxU41 ( 0 2679 ) COMPLEX( 390., 0.)
R_D52120xxU41 ( 2678 2666 )  100.n
R_D52120LOADxxU41 ( 0 2678 ) COMPLEX( 390., 0.)
R_D52121xxU41 ( 2677 2666 )  100.n
R_D52121LOADxxU41 ( 0 2677 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU41 ( 2676 2666 )  100.n
R_D52122LOADxxU41 ( 0 2676 ) COMPLEX( 151.656,-121.671)
R_D52123xxU41 ( 2675 2666 )  100.n
R_D52123LOADxxU41 ( 0 2675 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU41 ( 0 2673 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU41 ( 0 2674 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU41 ( 2674 2666 )  100.n
R_D52124xxU41 ( 2673 2666 )  100.n
R_D52125xxU41 ( 2672 2666 )  100.n
R_D52125LOADxxU41 ( 2672 0 ) COMPLEX( 390., 0.)
R_D52126xxU41 ( 2671 2666 )  100.n
R_D52126LOADxxU41 ( 2671 0 ) COMPLEX( 390., 0.)
R_D52127xxU41 ( 2670 2666 )  100.n
R_D52127LOADxxU41 ( 2670 0 ) COMPLEX( 390., 0.)
R_D52128xxU41 ( 2669 2666 )  100.n
R_D52128LOADxxU41 ( 2669 0 ) COMPLEX( 390., 0.)
R_D52129xxU41 ( 2668 2666 )  100.n
R_D52129LOADxxU41 ( 2668 0 ) COMPLEX( 390., 0.)
R_D52130xxU41 ( 2667 2666 )  100.n
R_D52130LOADxxU41 ( 2667 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU41 ( 2665 2666 )  100.n
R_D52131LOADxxU41 ( 2665 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U42CCM 
R_D52101xxU42 ( 2699 2730 )  100.n
R_D52101LOADxxU42 ( 0 2730 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU42 ( 2729 2699 )  100.n
R_D52102LOADxxU42 ( 0 2729 ) COMPLEX( 390., 0.)
R_D52103xxU42 ( 2728 2699 )  100.n
R_D52103LOADxxU42 ( 0 2728 ) COMPLEX( 390., 0.)
R_D52104xxU42 ( 2727 2699 )  100.n
R_D52104LOADxxU42 ( 0 2727 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU42 ( 2726 2699 )  100.n
R_D52105LOADxxU42 ( 0 2726 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU42 ( 2725 2699 )  100.n
R_D52106LOADxxU42 ( 0 2725 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU42 ( 0 2723 ) COMPLEX( 390., 0.)
R_D52108LOADxxU42 ( 0 2724 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU42 ( 2724 2699 )  100.n
R_D52107xxU42 ( 2723 2699 )  100.n
R_D52109xxU42 ( 2722 2699 )  100.n
R_D52109LOADxxU42 ( 2722 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU42 ( 2721 2699 )  100.n
R_D52110LOADxxU42 ( 2721 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU42 ( 2720 2699 )  100.n
R_D52111LOADxxU42 ( 2720 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU42 ( 2719 2699 )  100.n
R_D52112LOADxxU42 ( 2719 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU42 ( 2718 2699 )  100.n
R_D52113LOADxxU42 ( 2718 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU42 ( 2717 2699 )  100.n
R_D52114LOADxxU42 ( 2717 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU42 ( 2716 2699 )  100.n
R_D52116LOADxxU42 ( 2716 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU42 ( 538 2699 )  100.n
R_D52115xxU42 ( 2714 2699 )  100.n
R_D52115LOADxxU42 ( 2714 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU42 ( 2699 2713 )  100.n
R_D52118LOADxxU42 ( 0 2713 ) COMPLEX( 390., 0.)
R_D52119xxU42 ( 2712 2699 )  100.n
R_D52119LOADxxU42 ( 0 2712 ) COMPLEX( 390., 0.)
R_D52120xxU42 ( 2711 2699 )  100.n
R_D52120LOADxxU42 ( 0 2711 ) COMPLEX( 390., 0.)
R_D52121xxU42 ( 2710 2699 )  100.n
R_D52121LOADxxU42 ( 0 2710 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU42 ( 2709 2699 )  100.n
R_D52122LOADxxU42 ( 0 2709 ) COMPLEX( 151.656,-121.671)
R_D52123xxU42 ( 2708 2699 )  100.n
R_D52123LOADxxU42 ( 0 2708 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU42 ( 0 2706 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU42 ( 0 2707 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU42 ( 2707 2699 )  100.n
R_D52124xxU42 ( 2706 2699 )  100.n
R_D52125xxU42 ( 2705 2699 )  100.n
R_D52125LOADxxU42 ( 2705 0 ) COMPLEX( 390., 0.)
R_D52126xxU42 ( 2704 2699 )  100.n
R_D52126LOADxxU42 ( 2704 0 ) COMPLEX( 390., 0.)
R_D52127xxU42 ( 2703 2699 )  100.n
R_D52127LOADxxU42 ( 2703 0 ) COMPLEX( 390., 0.)
R_D52128xxU42 ( 2702 2699 )  100.n
R_D52128LOADxxU42 ( 2702 0 ) COMPLEX( 390., 0.)
R_D52129xxU42 ( 2701 2699 )  100.n
R_D52129LOADxxU42 ( 2701 0 ) COMPLEX( 390., 0.)
R_D52130xxU42 ( 2700 2699 )  100.n
R_D52130LOADxxU42 ( 2700 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU42 ( 2698 2699 )  100.n
R_D52131LOADxxU42 ( 2698 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U43CCM 
R_D52101xxU43 ( 2732 2763 )  100.n
R_D52101LOADxxU43 ( 0 2763 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU43 ( 2762 2732 )  100.n
R_D52102LOADxxU43 ( 0 2762 ) COMPLEX( 390., 0.)
R_D52103xxU43 ( 2761 2732 )  100.n
R_D52103LOADxxU43 ( 0 2761 ) COMPLEX( 390., 0.)
R_D52104xxU43 ( 2760 2732 )  100.n
R_D52104LOADxxU43 ( 0 2760 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU43 ( 2759 2732 )  100.n
R_D52105LOADxxU43 ( 0 2759 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU43 ( 2758 2732 )  100.n
R_D52106LOADxxU43 ( 0 2758 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU43 ( 0 2756 ) COMPLEX( 390., 0.)
R_D52108LOADxxU43 ( 0 2757 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU43 ( 2757 2732 )  100.n
R_D52107xxU43 ( 2756 2732 )  100.n
R_D52109xxU43 ( 2755 2732 )  100.n
R_D52109LOADxxU43 ( 2755 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU43 ( 2754 2732 )  100.n
R_D52110LOADxxU43 ( 2754 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU43 ( 2753 2732 )  100.n
R_D52111LOADxxU43 ( 2753 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU43 ( 2752 2732 )  100.n
R_D52112LOADxxU43 ( 2752 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU43 ( 2751 2732 )  100.n
R_D52113LOADxxU43 ( 2751 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU43 ( 2750 2732 )  100.n
R_D52114LOADxxU43 ( 2750 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU43 ( 2749 2732 )  100.n
R_D52116LOADxxU43 ( 2749 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU43 ( 539 2732 )  100.n
R_D52115xxU43 ( 2747 2732 )  100.n
R_D52115LOADxxU43 ( 2747 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU43 ( 2732 2746 )  100.n
R_D52118LOADxxU43 ( 0 2746 ) COMPLEX( 390., 0.)
R_D52119xxU43 ( 2745 2732 )  100.n
R_D52119LOADxxU43 ( 0 2745 ) COMPLEX( 390., 0.)
R_D52120xxU43 ( 2744 2732 )  100.n
R_D52120LOADxxU43 ( 0 2744 ) COMPLEX( 390., 0.)
R_D52121xxU43 ( 2743 2732 )  100.n
R_D52121LOADxxU43 ( 0 2743 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU43 ( 2742 2732 )  100.n
R_D52122LOADxxU43 ( 0 2742 ) COMPLEX( 151.656,-121.671)
R_D52123xxU43 ( 2741 2732 )  100.n
R_D52123LOADxxU43 ( 0 2741 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU43 ( 0 2739 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU43 ( 0 2740 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU43 ( 2740 2732 )  100.n
R_D52124xxU43 ( 2739 2732 )  100.n
R_D52125xxU43 ( 2738 2732 )  100.n
R_D52125LOADxxU43 ( 2738 0 ) COMPLEX( 390., 0.)
R_D52126xxU43 ( 2737 2732 )  100.n
R_D52126LOADxxU43 ( 2737 0 ) COMPLEX( 390., 0.)
R_D52127xxU43 ( 2736 2732 )  100.n
R_D52127LOADxxU43 ( 2736 0 ) COMPLEX( 390., 0.)
R_D52128xxU43 ( 2735 2732 )  100.n
R_D52128LOADxxU43 ( 2735 0 ) COMPLEX( 390., 0.)
R_D52129xxU43 ( 2734 2732 )  100.n
R_D52129LOADxxU43 ( 2734 0 ) COMPLEX( 390., 0.)
R_D52130xxU43 ( 2733 2732 )  100.n
R_D52130LOADxxU43 ( 2733 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU43 ( 2731 2732 )  100.n
R_D52131LOADxxU43 ( 2731 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U44CCM 
R_D52101xxU44 ( 2765 2796 )  100.n
R_D52101LOADxxU44 ( 0 2796 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU44 ( 2795 2765 )  100.n
R_D52102LOADxxU44 ( 0 2795 ) COMPLEX( 390., 0.)
R_D52103xxU44 ( 2794 2765 )  100.n
R_D52103LOADxxU44 ( 0 2794 ) COMPLEX( 390., 0.)
R_D52104xxU44 ( 2793 2765 )  100.n
R_D52104LOADxxU44 ( 0 2793 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU44 ( 2792 2765 )  100.n
R_D52105LOADxxU44 ( 0 2792 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU44 ( 2791 2765 )  100.n
R_D52106LOADxxU44 ( 0 2791 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU44 ( 0 2789 ) COMPLEX( 390., 0.)
R_D52108LOADxxU44 ( 0 2790 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU44 ( 2790 2765 )  100.n
R_D52107xxU44 ( 2789 2765 )  100.n
R_D52109xxU44 ( 2788 2765 )  100.n
R_D52109LOADxxU44 ( 2788 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU44 ( 2787 2765 )  100.n
R_D52110LOADxxU44 ( 2787 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU44 ( 2786 2765 )  100.n
R_D52111LOADxxU44 ( 2786 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU44 ( 2785 2765 )  100.n
R_D52112LOADxxU44 ( 2785 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU44 ( 2784 2765 )  100.n
R_D52113LOADxxU44 ( 2784 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU44 ( 2783 2765 )  100.n
R_D52114LOADxxU44 ( 2783 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU44 ( 2782 2765 )  100.n
R_D52116LOADxxU44 ( 2782 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU44 ( 542 2765 )  100.n
R_D52115xxU44 ( 2780 2765 )  100.n
R_D52115LOADxxU44 ( 2780 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU44 ( 2765 2779 )  100.n
R_D52118LOADxxU44 ( 0 2779 ) COMPLEX( 390., 0.)
R_D52119xxU44 ( 2778 2765 )  100.n
R_D52119LOADxxU44 ( 0 2778 ) COMPLEX( 390., 0.)
R_D52120xxU44 ( 2777 2765 )  100.n
R_D52120LOADxxU44 ( 0 2777 ) COMPLEX( 390., 0.)
R_D52121xxU44 ( 2776 2765 )  100.n
R_D52121LOADxxU44 ( 0 2776 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU44 ( 2775 2765 )  100.n
R_D52122LOADxxU44 ( 0 2775 ) COMPLEX( 151.656,-121.671)
R_D52123xxU44 ( 2774 2765 )  100.n
R_D52123LOADxxU44 ( 0 2774 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU44 ( 0 2772 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU44 ( 0 2773 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU44 ( 2773 2765 )  100.n
R_D52124xxU44 ( 2772 2765 )  100.n
R_D52125xxU44 ( 2771 2765 )  100.n
R_D52125LOADxxU44 ( 2771 0 ) COMPLEX( 390., 0.)
R_D52126xxU44 ( 2770 2765 )  100.n
R_D52126LOADxxU44 ( 2770 0 ) COMPLEX( 390., 0.)
R_D52127xxU44 ( 2769 2765 )  100.n
R_D52127LOADxxU44 ( 2769 0 ) COMPLEX( 390., 0.)
R_D52128xxU44 ( 2768 2765 )  100.n
R_D52128LOADxxU44 ( 2768 0 ) COMPLEX( 390., 0.)
R_D52129xxU44 ( 2767 2765 )  100.n
R_D52129LOADxxU44 ( 2767 0 ) COMPLEX( 390., 0.)
R_D52130xxU44 ( 2766 2765 )  100.n
R_D52130LOADxxU44 ( 2766 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU44 ( 2764 2765 )  100.n
R_D52131LOADxxU44 ( 2764 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U45CCM 
R_D52101xxU45 ( 2798 2829 )  100.n
R_D52101LOADxxU45 ( 0 2829 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU45 ( 2828 2798 )  100.n
R_D52102LOADxxU45 ( 0 2828 ) COMPLEX( 390., 0.)
R_D52103xxU45 ( 2827 2798 )  100.n
R_D52103LOADxxU45 ( 0 2827 ) COMPLEX( 390., 0.)
R_D52104xxU45 ( 2826 2798 )  100.n
R_D52104LOADxxU45 ( 0 2826 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU45 ( 2825 2798 )  100.n
R_D52105LOADxxU45 ( 0 2825 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU45 ( 2824 2798 )  100.n
R_D52106LOADxxU45 ( 0 2824 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU45 ( 0 2822 ) COMPLEX( 390., 0.)
R_D52108LOADxxU45 ( 0 2823 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU45 ( 2823 2798 )  100.n
R_D52107xxU45 ( 2822 2798 )  100.n
R_D52109xxU45 ( 2821 2798 )  100.n
R_D52109LOADxxU45 ( 2821 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU45 ( 2820 2798 )  100.n
R_D52110LOADxxU45 ( 2820 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU45 ( 2819 2798 )  100.n
R_D52111LOADxxU45 ( 2819 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU45 ( 2818 2798 )  100.n
R_D52112LOADxxU45 ( 2818 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU45 ( 2817 2798 )  100.n
R_D52113LOADxxU45 ( 2817 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU45 ( 2816 2798 )  100.n
R_D52114LOADxxU45 ( 2816 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU45 ( 2815 2798 )  100.n
R_D52116LOADxxU45 ( 2815 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU45 ( 411 2798 )  100.n
R_D52115xxU45 ( 2813 2798 )  100.n
R_D52115LOADxxU45 ( 2813 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU45 ( 2798 2812 )  100.n
R_D52118LOADxxU45 ( 0 2812 ) COMPLEX( 390., 0.)
R_D52119xxU45 ( 2811 2798 )  100.n
R_D52119LOADxxU45 ( 0 2811 ) COMPLEX( 390., 0.)
R_D52120xxU45 ( 2810 2798 )  100.n
R_D52120LOADxxU45 ( 0 2810 ) COMPLEX( 390., 0.)
R_D52121xxU45 ( 2809 2798 )  100.n
R_D52121LOADxxU45 ( 0 2809 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU45 ( 2808 2798 )  100.n
R_D52122LOADxxU45 ( 0 2808 ) COMPLEX( 151.656,-121.671)
R_D52123xxU45 ( 2807 2798 )  100.n
R_D52123LOADxxU45 ( 0 2807 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU45 ( 0 2805 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU45 ( 0 2806 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU45 ( 2806 2798 )  100.n
R_D52124xxU45 ( 2805 2798 )  100.n
R_D52125xxU45 ( 2804 2798 )  100.n
R_D52125LOADxxU45 ( 2804 0 ) COMPLEX( 390., 0.)
R_D52126xxU45 ( 2803 2798 )  100.n
R_D52126LOADxxU45 ( 2803 0 ) COMPLEX( 390., 0.)
R_D52127xxU45 ( 2802 2798 )  100.n
R_D52127LOADxxU45 ( 2802 0 ) COMPLEX( 390., 0.)
R_D52128xxU45 ( 2801 2798 )  100.n
R_D52128LOADxxU45 ( 2801 0 ) COMPLEX( 390., 0.)
R_D52129xxU45 ( 2800 2798 )  100.n
R_D52129LOADxxU45 ( 2800 0 ) COMPLEX( 390., 0.)
R_D52130xxU45 ( 2799 2798 )  100.n
R_D52130LOADxxU45 ( 2799 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU45 ( 2797 2798 )  100.n
R_D52131LOADxxU45 ( 2797 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U46CCM 
R_D52101xxU46 ( 2831 2862 )  100.n
R_D52101LOADxxU46 ( 0 2862 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU46 ( 2861 2831 )  100.n
R_D52102LOADxxU46 ( 0 2861 ) COMPLEX( 390., 0.)
R_D52103xxU46 ( 2860 2831 )  100.n
R_D52103LOADxxU46 ( 0 2860 ) COMPLEX( 390., 0.)
R_D52104xxU46 ( 2859 2831 )  100.n
R_D52104LOADxxU46 ( 0 2859 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU46 ( 2858 2831 )  100.n
R_D52105LOADxxU46 ( 0 2858 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU46 ( 2857 2831 )  100.n
R_D52106LOADxxU46 ( 0 2857 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU46 ( 0 2855 ) COMPLEX( 390., 0.)
R_D52108LOADxxU46 ( 0 2856 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU46 ( 2856 2831 )  100.n
R_D52107xxU46 ( 2855 2831 )  100.n
R_D52109xxU46 ( 2854 2831 )  100.n
R_D52109LOADxxU46 ( 2854 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU46 ( 2853 2831 )  100.n
R_D52110LOADxxU46 ( 2853 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU46 ( 2852 2831 )  100.n
R_D52111LOADxxU46 ( 2852 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU46 ( 2851 2831 )  100.n
R_D52112LOADxxU46 ( 2851 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU46 ( 2850 2831 )  100.n
R_D52113LOADxxU46 ( 2850 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU46 ( 2849 2831 )  100.n
R_D52114LOADxxU46 ( 2849 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU46 ( 2848 2831 )  100.n
R_D52116LOADxxU46 ( 2848 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU46 ( 413 2831 )  100.n
R_D52115xxU46 ( 2846 2831 )  100.n
R_D52115LOADxxU46 ( 2846 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU46 ( 2831 2845 )  100.n
R_D52118LOADxxU46 ( 0 2845 ) COMPLEX( 390., 0.)
R_D52119xxU46 ( 2844 2831 )  100.n
R_D52119LOADxxU46 ( 0 2844 ) COMPLEX( 390., 0.)
R_D52120xxU46 ( 2843 2831 )  100.n
R_D52120LOADxxU46 ( 0 2843 ) COMPLEX( 390., 0.)
R_D52121xxU46 ( 2842 2831 )  100.n
R_D52121LOADxxU46 ( 0 2842 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU46 ( 2841 2831 )  100.n
R_D52122LOADxxU46 ( 0 2841 ) COMPLEX( 151.656,-121.671)
R_D52123xxU46 ( 2840 2831 )  100.n
R_D52123LOADxxU46 ( 0 2840 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU46 ( 0 2838 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU46 ( 0 2839 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU46 ( 2839 2831 )  100.n
R_D52124xxU46 ( 2838 2831 )  100.n
R_D52125xxU46 ( 2837 2831 )  100.n
R_D52125LOADxxU46 ( 2837 0 ) COMPLEX( 390., 0.)
R_D52126xxU46 ( 2836 2831 )  100.n
R_D52126LOADxxU46 ( 2836 0 ) COMPLEX( 390., 0.)
R_D52127xxU46 ( 2835 2831 )  100.n
R_D52127LOADxxU46 ( 2835 0 ) COMPLEX( 390., 0.)
R_D52128xxU46 ( 2834 2831 )  100.n
R_D52128LOADxxU46 ( 2834 0 ) COMPLEX( 390., 0.)
R_D52129xxU46 ( 2833 2831 )  100.n
R_D52129LOADxxU46 ( 2833 0 ) COMPLEX( 390., 0.)
R_D52130xxU46 ( 2832 2831 )  100.n
R_D52130LOADxxU46 ( 2832 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU46 ( 2830 2831 )  100.n
R_D52131LOADxxU46 ( 2830 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U47CCM 
R_D52101xxU47 ( 2864 2895 )  100.n
R_D52101LOADxxU47 ( 0 2895 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU47 ( 2894 2864 )  100.n
R_D52102LOADxxU47 ( 0 2894 ) COMPLEX( 390., 0.)
R_D52103xxU47 ( 2893 2864 )  100.n
R_D52103LOADxxU47 ( 0 2893 ) COMPLEX( 390., 0.)
R_D52104xxU47 ( 2892 2864 )  100.n
R_D52104LOADxxU47 ( 0 2892 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU47 ( 2891 2864 )  100.n
R_D52105LOADxxU47 ( 0 2891 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU47 ( 2890 2864 )  100.n
R_D52106LOADxxU47 ( 0 2890 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU47 ( 0 2888 ) COMPLEX( 390., 0.)
R_D52108LOADxxU47 ( 0 2889 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU47 ( 2889 2864 )  100.n
R_D52107xxU47 ( 2888 2864 )  100.n
R_D52109xxU47 ( 2887 2864 )  100.n
R_D52109LOADxxU47 ( 2887 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU47 ( 2886 2864 )  100.n
R_D52110LOADxxU47 ( 2886 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU47 ( 2885 2864 )  100.n
R_D52111LOADxxU47 ( 2885 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU47 ( 2884 2864 )  100.n
R_D52112LOADxxU47 ( 2884 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU47 ( 2883 2864 )  100.n
R_D52113LOADxxU47 ( 2883 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU47 ( 2882 2864 )  100.n
R_D52114LOADxxU47 ( 2882 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU47 ( 2881 2864 )  100.n
R_D52116LOADxxU47 ( 2881 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU47 ( 417 2864 )  100.n
R_D52115xxU47 ( 2879 2864 )  100.n
R_D52115LOADxxU47 ( 2879 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU47 ( 2864 2878 )  100.n
R_D52118LOADxxU47 ( 0 2878 ) COMPLEX( 390., 0.)
R_D52119xxU47 ( 2877 2864 )  100.n
R_D52119LOADxxU47 ( 0 2877 ) COMPLEX( 390., 0.)
R_D52120xxU47 ( 2876 2864 )  100.n
R_D52120LOADxxU47 ( 0 2876 ) COMPLEX( 390., 0.)
R_D52121xxU47 ( 2875 2864 )  100.n
R_D52121LOADxxU47 ( 0 2875 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU47 ( 2874 2864 )  100.n
R_D52122LOADxxU47 ( 0 2874 ) COMPLEX( 151.656,-121.671)
R_D52123xxU47 ( 2873 2864 )  100.n
R_D52123LOADxxU47 ( 0 2873 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU47 ( 0 2871 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU47 ( 0 2872 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU47 ( 2872 2864 )  100.n
R_D52124xxU47 ( 2871 2864 )  100.n
R_D52125xxU47 ( 2870 2864 )  100.n
R_D52125LOADxxU47 ( 2870 0 ) COMPLEX( 390., 0.)
R_D52126xxU47 ( 2869 2864 )  100.n
R_D52126LOADxxU47 ( 2869 0 ) COMPLEX( 390., 0.)
R_D52127xxU47 ( 2868 2864 )  100.n
R_D52127LOADxxU47 ( 2868 0 ) COMPLEX( 390., 0.)
R_D52128xxU47 ( 2867 2864 )  100.n
R_D52128LOADxxU47 ( 2867 0 ) COMPLEX( 390., 0.)
R_D52129xxU47 ( 2866 2864 )  100.n
R_D52129LOADxxU47 ( 2866 0 ) COMPLEX( 390., 0.)
R_D52130xxU47 ( 2865 2864 )  100.n
R_D52130LOADxxU47 ( 2865 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU47 ( 2863 2864 )  100.n
R_D52131LOADxxU47 ( 2863 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U48CCM 
R_D52101xxU48 ( 2897 2928 )  100.n
R_D52101LOADxxU48 ( 0 2928 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU48 ( 2927 2897 )  100.n
R_D52102LOADxxU48 ( 0 2927 ) COMPLEX( 390., 0.)
R_D52103xxU48 ( 2926 2897 )  100.n
R_D52103LOADxxU48 ( 0 2926 ) COMPLEX( 390., 0.)
R_D52104xxU48 ( 2925 2897 )  100.n
R_D52104LOADxxU48 ( 0 2925 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU48 ( 2924 2897 )  100.n
R_D52105LOADxxU48 ( 0 2924 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU48 ( 2923 2897 )  100.n
R_D52106LOADxxU48 ( 0 2923 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU48 ( 0 2921 ) COMPLEX( 390., 0.)
R_D52108LOADxxU48 ( 0 2922 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU48 ( 2922 2897 )  100.n
R_D52107xxU48 ( 2921 2897 )  100.n
R_D52109xxU48 ( 2920 2897 )  100.n
R_D52109LOADxxU48 ( 2920 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU48 ( 2919 2897 )  100.n
R_D52110LOADxxU48 ( 2919 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU48 ( 2918 2897 )  100.n
R_D52111LOADxxU48 ( 2918 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU48 ( 2917 2897 )  100.n
R_D52112LOADxxU48 ( 2917 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU48 ( 2916 2897 )  100.n
R_D52113LOADxxU48 ( 2916 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU48 ( 2915 2897 )  100.n
R_D52114LOADxxU48 ( 2915 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU48 ( 2914 2897 )  100.n
R_D52116LOADxxU48 ( 2914 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU48 ( 416 2897 )  100.n
R_D52115xxU48 ( 2912 2897 )  100.n
R_D52115LOADxxU48 ( 2912 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU48 ( 2897 2911 )  100.n
R_D52118LOADxxU48 ( 0 2911 ) COMPLEX( 390., 0.)
R_D52119xxU48 ( 2910 2897 )  100.n
R_D52119LOADxxU48 ( 0 2910 ) COMPLEX( 390., 0.)
R_D52120xxU48 ( 2909 2897 )  100.n
R_D52120LOADxxU48 ( 0 2909 ) COMPLEX( 390., 0.)
R_D52121xxU48 ( 2908 2897 )  100.n
R_D52121LOADxxU48 ( 0 2908 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU48 ( 2907 2897 )  100.n
R_D52122LOADxxU48 ( 0 2907 ) COMPLEX( 151.656,-121.671)
R_D52123xxU48 ( 2906 2897 )  100.n
R_D52123LOADxxU48 ( 0 2906 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU48 ( 0 2904 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU48 ( 0 2905 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU48 ( 2905 2897 )  100.n
R_D52124xxU48 ( 2904 2897 )  100.n
R_D52125xxU48 ( 2903 2897 )  100.n
R_D52125LOADxxU48 ( 2903 0 ) COMPLEX( 390., 0.)
R_D52126xxU48 ( 2902 2897 )  100.n
R_D52126LOADxxU48 ( 2902 0 ) COMPLEX( 390., 0.)
R_D52127xxU48 ( 2901 2897 )  100.n
R_D52127LOADxxU48 ( 2901 0 ) COMPLEX( 390., 0.)
R_D52128xxU48 ( 2900 2897 )  100.n
R_D52128LOADxxU48 ( 2900 0 ) COMPLEX( 390., 0.)
R_D52129xxU48 ( 2899 2897 )  100.n
R_D52129LOADxxU48 ( 2899 0 ) COMPLEX( 390., 0.)
R_D52130xxU48 ( 2898 2897 )  100.n
R_D52130LOADxxU48 ( 2898 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU48 ( 2896 2897 )  100.n
R_D52131LOADxxU48 ( 2896 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U49CCM 
R_D52101xxU49 ( 2930 2961 )  100.n
R_D52101LOADxxU49 ( 0 2961 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU49 ( 2960 2930 )  100.n
R_D52102LOADxxU49 ( 0 2960 ) COMPLEX( 390., 0.)
R_D52103xxU49 ( 2959 2930 )  100.n
R_D52103LOADxxU49 ( 0 2959 ) COMPLEX( 390., 0.)
R_D52104xxU49 ( 2958 2930 )  100.n
R_D52104LOADxxU49 ( 0 2958 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU49 ( 2957 2930 )  100.n
R_D52105LOADxxU49 ( 0 2957 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU49 ( 2956 2930 )  100.n
R_D52106LOADxxU49 ( 0 2956 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU49 ( 0 2954 ) COMPLEX( 390., 0.)
R_D52108LOADxxU49 ( 0 2955 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU49 ( 2955 2930 )  100.n
R_D52107xxU49 ( 2954 2930 )  100.n
R_D52109xxU49 ( 2953 2930 )  100.n
R_D52109LOADxxU49 ( 2953 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU49 ( 2952 2930 )  100.n
R_D52110LOADxxU49 ( 2952 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU49 ( 2951 2930 )  100.n
R_D52111LOADxxU49 ( 2951 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU49 ( 2950 2930 )  100.n
R_D52112LOADxxU49 ( 2950 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU49 ( 2949 2930 )  100.n
R_D52113LOADxxU49 ( 2949 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU49 ( 2948 2930 )  100.n
R_D52114LOADxxU49 ( 2948 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU49 ( 2947 2930 )  100.n
R_D52116LOADxxU49 ( 2947 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU49 ( 399 2930 )  100.n
R_D52115xxU49 ( 2945 2930 )  100.n
R_D52115LOADxxU49 ( 2945 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU49 ( 2930 2944 )  100.n
R_D52118LOADxxU49 ( 0 2944 ) COMPLEX( 390., 0.)
R_D52119xxU49 ( 2943 2930 )  100.n
R_D52119LOADxxU49 ( 0 2943 ) COMPLEX( 390., 0.)
R_D52120xxU49 ( 2942 2930 )  100.n
R_D52120LOADxxU49 ( 0 2942 ) COMPLEX( 390., 0.)
R_D52121xxU49 ( 2941 2930 )  100.n
R_D52121LOADxxU49 ( 0 2941 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU49 ( 2940 2930 )  100.n
R_D52122LOADxxU49 ( 0 2940 ) COMPLEX( 151.656,-121.671)
R_D52123xxU49 ( 2939 2930 )  100.n
R_D52123LOADxxU49 ( 0 2939 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU49 ( 0 2937 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU49 ( 0 2938 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU49 ( 2938 2930 )  100.n
R_D52124xxU49 ( 2937 2930 )  100.n
R_D52125xxU49 ( 2936 2930 )  100.n
R_D52125LOADxxU49 ( 2936 0 ) COMPLEX( 390., 0.)
R_D52126xxU49 ( 2935 2930 )  100.n
R_D52126LOADxxU49 ( 2935 0 ) COMPLEX( 390., 0.)
R_D52127xxU49 ( 2934 2930 )  100.n
R_D52127LOADxxU49 ( 2934 0 ) COMPLEX( 390., 0.)
R_D52128xxU49 ( 2933 2930 )  100.n
R_D52128LOADxxU49 ( 2933 0 ) COMPLEX( 390., 0.)
R_D52129xxU49 ( 2932 2930 )  100.n
R_D52129LOADxxU49 ( 2932 0 ) COMPLEX( 390., 0.)
R_D52130xxU49 ( 2931 2930 )  100.n
R_D52130LOADxxU49 ( 2931 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU49 ( 2929 2930 )  100.n
R_D52131LOADxxU49 ( 2929 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA U50CCM 
R_D52101xxU50 ( 2963 2994 )  100.n
R_D52101LOADxxU50 ( 0 2994 ) COMPLEX( 1.4892,-0.8037)
R_D52102xxU50 ( 2993 2963 )  100.n
R_D52102LOADxxU50 ( 0 2993 ) COMPLEX( 390., 0.)
R_D52103xxU50 ( 2992 2963 )  100.n
R_D52103LOADxxU50 ( 0 2992 ) COMPLEX( 390., 0.)
R_D52104xxU50 ( 2991 2963 )  100.n
R_D52104LOADxxU50 ( 0 2991 ) COMPLEX( 517.44,-527.8944)
R_D52105xxU50 ( 2990 2963 )  100.n
R_D52105LOADxxU50 ( 0 2990 ) COMPLEX( 11.6097,-6.8889)
R_D52106xxU50 ( 2989 2963 )  100.n
R_D52106LOADxxU50 ( 0 2989 ) COMPLEX( 11.6097,-6.8889)
R_D52107LOADxxU50 ( 0 2987 ) COMPLEX( 390., 0.)
R_D52108LOADxxU50 ( 0 2988 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxU50 ( 2988 2963 )  100.n
R_D52107xxU50 ( 2987 2963 )  100.n
R_D52109xxU50 ( 2986 2963 )  100.n
R_D52109LOADxxU50 ( 2986 0 ) COMPLEX( 9.7692,-5.5365)
R_D52110xxU50 ( 2985 2963 )  100.n
R_D52110LOADxxU50 ( 2985 0 ) COMPLEX( 168.96,-126.72)
R_D52111xxU50 ( 2984 2963 )  100.n
R_D52111LOADxxU50 ( 2984 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxU50 ( 2983 2963 )  100.n
R_D52112LOADxxU50 ( 2983 0 ) COMPLEX( 3.1791,-1.9701)
R_D52113xxU50 ( 2982 2963 )  100.n
R_D52113LOADxxU50 ( 2982 0 ) COMPLEX( 3.1791,-1.9701)
R_D52114xxU50 ( 2981 2963 )  100.n
R_D52114LOADxxU50 ( 2981 0 ) COMPLEX( 168.96,-126.72)
R_D52116xxU50 ( 2980 2963 )  100.n
R_D52116LOADxxU50 ( 2980 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52ExxU50 ( 404 2963 )  100.n
R_D52115xxU50 ( 2978 2963 )  100.n
R_D52115LOADxxU50 ( 2978 0 ) COMPLEX( 1.363267K,-1.593835K)
R_D52118xxU50 ( 2963 2977 )  100.n
R_D52118LOADxxU50 ( 0 2977 ) COMPLEX( 390., 0.)
R_D52119xxU50 ( 2976 2963 )  100.n
R_D52119LOADxxU50 ( 0 2976 ) COMPLEX( 390., 0.)
R_D52120xxU50 ( 2975 2963 )  100.n
R_D52120LOADxxU50 ( 0 2975 ) COMPLEX( 390., 0.)
R_D52121xxU50 ( 2974 2963 )  100.n
R_D52121LOADxxU50 ( 0 2974 ) COMPLEX( 26.6742,-17.9253)
R_D52122xxU50 ( 2973 2963 )  100.n
R_D52122LOADxxU50 ( 0 2973 ) COMPLEX( 151.656,-121.671)
R_D52123xxU50 ( 2972 2963 )  100.n
R_D52123LOADxxU50 ( 0 2972 ) COMPLEX( 168.96,-126.72)
R_D52124LOADxxU50 ( 0 2970 ) COMPLEX( 168.96,-126.72)
R_D52117LOADxxU50 ( 0 2971 ) COMPLEX( 1.363267K,-1.593835K)
R_D52117xxU50 ( 2971 2963 )  100.n
R_D52124xxU50 ( 2970 2963 )  100.n
R_D52125xxU50 ( 0 0 )  1.E+12
R_D52125LOADxxU50 ( 2969 0 ) COMPLEX( 390., 0.)
R_D52126xxU50 ( 2968 2963 )  100.n
R_D52126LOADxxU50 ( 2968 0 ) COMPLEX( 390., 0.)
R_D52127xxU50 ( 2967 2963 )  100.n
R_D52127LOADxxU50 ( 2967 0 ) COMPLEX( 390., 0.)
R_D52128xxU50 ( 2966 2963 )  100.n
R_D52128LOADxxU50 ( 2966 0 ) COMPLEX( 390., 0.)
R_D52129xxU50 ( 0 0 )  1.E+12
R_D52129LOADxxU50 ( 2965 0 ) COMPLEX( 390., 0.)
R_D52130xxU50 ( 2964 2963 )  100.n
R_D52130LOADxxU50 ( 2964 0 ) COMPLEX( 168.96,-126.72)
R_D52131xxU50 ( 2962 2963 )  100.n
R_D52131LOADxxU50 ( 2962 0 ) COMPLEX( 168.96,-126.72)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG8 
R_D52101xxQSG8 ( 2996 3062 )  100.n
R_D52101LOADxxQSG8 ( 0 3062 ) COMPLEX( 53.3484,-35.8503)
R_D52102xxQSG8 ( 3061 2996 )  100.n
R_D52102LOADxxQSG8 ( 0 3061 ) COMPLEX( 390., 0.)
R_D52103xxQSG8 ( 3060 2996 )  100.n
R_D52103LOADxxQSG8 ( 0 3060 ) COMPLEX( 86.7843,-60.576)
R_D52104xxQSG8 ( 3059 2996 )  100.n
R_D52104LOADxxQSG8 ( 0 3059 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG8 ( 3058 2996 )  100.n
R_D52105LOADxxQSG8 ( 0 3058 ) COMPLEX( 3.9963,-2.265)
R_D52106xxQSG8 ( 3057 2996 )  100.n
R_D52106LOADxxQSG8 ( 0 3057 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG8 ( 0 3056 ) COMPLEX( 390., 0.)
R_D52108xxQSG8 ( 3056 2996 )  100.n
R_D52112xxQSG8 ( 3055 2996 )  100.n
R_D52112LOADxxQSG8 ( 3055 0 ) COMPLEX( 102.99,-74.5635)
R_D52113xxQSG8 ( 3054 2996 )  100.n
R_D52113LOADxxQSG8 ( 3054 0 ) COMPLEX( 418.2288,-214.2651)
R_D52114xxQSG8 ( 3053 2996 )  100.n
R_D52114LOADxxQSG8 ( 3053 0 ) COMPLEX( 3.9963,-2.265)
R_D52115xxQSG8 ( 3052 2996 )  100.n
R_D52115LOADxxQSG8 ( 3052 0 ) COMPLEX( 390., 0.)
R_D52116xxQSG8 ( 3051 2996 )  100.n
R_D52116LOADxxQSG8 ( 3051 0 ) COMPLEX( 390., 0.)
R_D52117xxQSG8 ( 3050 2996 )  100.n
R_D52117LOADxxQSG8 ( 3050 0 ) COMPLEX( 13.9875,-8.6688)
R_D52L1xxQSG8 ( 0 0 )  1.E+12
R_D52118xxQSG8 ( 3048 2996 )  100.n
R_D52118LOADxxQSG8 ( 3048 0 ) COMPLEX( 30.976, 0.)
R_D52111xxQSG8 ( 3047 2996 )  100.n
R_D52111LOADxxQSG8 ( 3047 0 ) COMPLEX( 390., 0.)
R_D52119xxQSG8 ( 3046 2996 )  100.n
R_D52119LOADxxQSG8 ( 3046 0 ) COMPLEX( 8.1777,-4.4139)
R_D52120xxQSG8 ( 3045 2996 )  100.n
R_D52120LOADxxQSG8 ( 3045 0 ) COMPLEX( 3.9963,-2.265)
R_D52109LOADxxQSG8 ( 0 3044 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG8 ( 3044 2996 )  100.n
R_D52107LOADxxQSG8 ( 0 0 )  1.E+12
R_D52107xxQSG8 ( 3043 2996 )  100.n
R_D52L2xxQSG8 ( 2998 3023 )  100.n
R_D52E2xxQSG8 ( 481 3023 )  100.n
R_D52E1xxQSG8 ( 603 2996 )  100.n
R_D52201xxQSG8 ( 3023 3040 )  100.n
R_D52201LOADxxQSG8 ( 0 3040 ) COMPLEX( 42.4488,-29.6295)
R_D52202xxQSG8 ( 3039 3023 )  100.n
R_D52202LOADxxQSG8 ( 0 3039 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG8 ( 3038 3023 )  100.n
R_D52203LOADxxQSG8 ( 0 3038 ) COMPLEX( 390., 0.)
R_D52204xxQSG8 ( 3037 3023 )  100.n
R_D52204LOADxxQSG8 ( 0 3037 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG8 ( 3036 3023 )  100.n
R_D52205LOADxxQSG8 ( 0 3036 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG8 ( 3035 3023 )  100.n
R_D52206LOADxxQSG8 ( 0 0 )  1.E+12
R_D52208LOADxxQSG8 ( 0 3034 ) COMPLEX( 235.5726,-188.9955)
R_D52208xxQSG8 ( 3034 3023 )  100.n
R_D52211xxQSG8 ( 3033 3023 )  100.n
R_D52211LOADxxQSG8 ( 3033 0 ) COMPLEX( 235.5726,-188.9955)
R_D52212xxQSG8 ( 3032 3023 )  100.n
R_D52212LOADxxQSG8 ( 3032 0 ) COMPLEX( 390., 0.)
R_D52213xxQSG8 ( 3031 3023 )  100.n
R_D52213LOADxxQSG8 ( 3031 0 ) COMPLEX( 418.2288,-214.2651)
R_D52214xxQSG8 ( 3030 3023 )  100.n
R_D52214LOADxxQSG8 ( 3030 0 ) COMPLEX( 13.9875,-8.6688)
R_D52215xxQSG8 ( 3029 3023 )  100.n
R_D52215LOADxxQSG8 ( 3029 0 ) COMPLEX( 390., 0.)
R_D52216xxQSG8 ( 3028 3023 )  100.n
R_D52216LOADxxQSG8 ( 3028 0 ) COMPLEX( 8.1777,-4.4139)
R_D52217xxQSG8 ( 3027 3023 )  100.n
R_D52217LOADxxQSG8 ( 3027 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG8 ( 3026 3023 )  100.n
R_D52210LOADxxQSG8 ( 3026 0 ) COMPLEX( 390., 0.)
R_D52218xxQSG8 ( 3025 3023 )  100.n
R_D52218LOADxxQSG8 ( 3025 0 ) COMPLEX( 3.9963,-2.265)
R_D52209LOADxxQSG8 ( 0 3024 ) COMPLEX( 3.9963,-2.265)
R_D52209xxQSG8 ( 3024 3023 )  100.n
R_D52207LOADxxQSG8 ( 3022 0 ) COMPLEX( 418.2288,-214.2651)
R_D52207xxQSG8 ( 3022 3023 )  100.n
R_D52301xxQSG8 ( 2998 3020 )  100.n
R_D52301LOADxxQSG8 ( 0 3020 ) COMPLEX( 2.0445,-1.1034)
R_D52302xxQSG8 ( 3019 2998 )  100.n
R_D52302LOADxxQSG8 ( 0 3019 ) COMPLEX( 390., 0.)
R_D52303xxQSG8 ( 3018 2998 )  100.n
R_D52303LOADxxQSG8 ( 0 3018 ) COMPLEX( 176.6793,-141.7467)
R_D52304xxQSG8 ( 3017 2998 )  100.n
R_D52304LOADxxQSG8 ( 0 3017 ) COMPLEX( 21.6276,-14.5338)
R_D52305xxQSG8 ( 3016 2998 )  100.n
R_D52305LOADxxQSG8 ( 0 3016 ) COMPLEX( 390., 0.)
R_D52306xxQSG8 ( 3015 2998 )  100.n
R_D52306LOADxxQSG8 ( 0 3015 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG8 ( 0 3014 ) COMPLEX( 86.7843,-60.576)
R_D52308xxQSG8 ( 3014 2998 )  100.n
R_D52311xxQSG8 ( 3013 2998 )  100.n
R_D52311LOADxxQSG8 ( 3013 0 ) COMPLEX( 390., 0.)
R_D52312xxQSG8 ( 3012 2998 )  100.n
R_D52312LOADxxQSG8 ( 3012 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG8 ( 3011 2998 )  100.n
R_D52313LOADxxQSG8 ( 3011 0 ) COMPLEX( 168.96,-126.72)
R_D52314xxQSG8 ( 3010 2998 )  100.n
R_D52314LOADxxQSG8 ( 3010 0 ) COMPLEX( 390., 0.)
R_D52315xxQSG8 ( 3009 2998 )  100.n
R_D52315LOADxxQSG8 ( 3009 0 ) COMPLEX( 2.4495,-0.8052)
R_D52316xxQSG8 ( 3008 2998 )  100.n
R_D52316LOADxxQSG8 ( 3008 0 ) COMPLEX( 168.96,-126.72)
R_D52317xxQSG8 ( 3007 2998 )  100.n
R_D52317LOADxxQSG8 ( 3007 0 ) COMPLEX( 6.078,-3.2805)
R_D52310xxQSG8 ( 3006 2998 )  100.n
R_D52310LOADxxQSG8 ( 3006 0 ) COMPLEX( 390., 0.)
R_D52318xxQSG8 ( 3005 2998 )  100.n
R_D52318LOADxxQSG8 ( 3005 0 ) COMPLEX( 6.078,-3.2805)
R_D52319xxQSG8 ( 3004 2998 )  100.n
R_D52319LOADxxQSG8 ( 3004 0 ) COMPLEX( 6.078,-3.2805)
R_D52309LOADxxQSG8 ( 0 3003 ) COMPLEX( 390., 0.)
R_D52309xxQSG8 ( 3003 2998 )  100.n
R_D52307LOADxxQSG8 ( 3002 0 ) COMPLEX( 390., 0.)
R_D52307xxQSG8 ( 3002 2998 )  100.n
R_D52320xxQSG8 ( 2998 3001 )  100.n
R_D52320LOADxxQSG8 ( 0 3001 ) COMPLEX( 10.7391,-6.372)
R_D52321xxQSG8 ( 3000 2998 )  100.n
R_D52321LOADxxQSG8 ( 0 3000 ) COMPLEX( 10.7391,-6.372)
R_D52323xxQSG8 ( 2999 2998 )  100.n
R_D52323LOADxxQSG8 ( 2999 0 ) COMPLEX( 2.4495,-0.8052)
R_D52322xxQSG8 ( 2997 2998 )  100.n
R_D52322LOADxxQSG8 ( 2997 0 ) COMPLEX( 390., 0.)
R_D52110LOADxxQSG8 ( 0 2995 ) COMPLEX( 3.9963,-2.265)
R_D52110xxQSG8 ( 2995 2996 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG9 
R_D52101xxQSG9 ( 3064 3114 )  100.n
R_D52101LOADxxQSG9 ( 0 3114 ) COMPLEX( 390., 0.)
R_D52102xxQSG9 ( 3113 3064 )  100.n
R_D52102LOADxxQSG9 ( 0 3113 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG9 ( 3112 3064 )  100.n
R_D52103LOADxxQSG9 ( 0 3112 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG9 ( 3111 3064 )  100.n
R_D52104LOADxxQSG9 ( 0 3111 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG9 ( 3110 3064 )  100.n
R_D52105LOADxxQSG9 ( 0 3110 ) COMPLEX( 30.976, 0.)
R_D52106xxQSG9 ( 3109 3064 )  100.n
R_D52106LOADxxQSG9 ( 0 0 )  1.E+12
R_D52108LOADxxQSG9 ( 0 3108 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG9 ( 3108 3064 )  100.n
R_D52111xxQSG9 ( 3107 3064 )  100.n
R_D52111LOADxxQSG9 ( 3107 0 ) COMPLEX( 8.1777,-4.4139)
R_D52112xxQSG9 ( 3106 3064 )  100.n
R_D52112LOADxxQSG9 ( 3106 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG9 ( 3105 3064 )  100.n
R_D52113LOADxxQSG9 ( 3105 0 ) COMPLEX( 390., 0.)
R_D52L1xxQSG9 ( 0 0 )  1.E+12
R_D52110xxQSG9 ( 3103 3064 )  100.n
R_D52110LOADxxQSG9 ( 3103 0 ) COMPLEX( 418.2288,-214.2651)
R_D52109LOADxxQSG9 ( 0 3102 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG9 ( 3102 3064 )  100.n
R_D52107LOADxxQSG9 ( 3101 0 ) COMPLEX( 10.7391,-6.372)
R_D52107xxQSG9 ( 3101 3064 )  100.n
R_D52L2xxQSG9 ( 3082 3067 )  100.n
R_D52E2xxQSG9 ( 608 3067 )  100.n
R_D52E1xxQSG9 ( 487 3064 )  100.n
R_D52301xxQSG9 ( 3082 3098 )  100.n
R_D52301LOADxxQSG9 ( 0 3098 ) COMPLEX( 1.9074,-1.182)
R_D52302xxQSG9 ( 3097 3082 )  100.n
R_D52302LOADxxQSG9 ( 0 3097 ) COMPLEX( 390., 0.)
R_D52303xxQSG9 ( 3096 3082 )  100.n
R_D52303LOADxxQSG9 ( 0 3096 ) COMPLEX( 390., 0.)
R_D52304xxQSG9 ( 3095 3082 )  100.n
R_D52304LOADxxQSG9 ( 0 3095 ) COMPLEX( 390., 0.)
R_D52305xxQSG9 ( 3094 3082 )  100.n
R_D52305LOADxxQSG9 ( 0 3094 ) COMPLEX( 390., 0.)
R_D52306xxQSG9 ( 3093 3082 )  100.n
R_D52306LOADxxQSG9 ( 0 3093 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG9 ( 0 3092 ) COMPLEX( 390., 0.)
R_D52308xxQSG9 ( 3092 3082 )  100.n
R_D52311xxQSG9 ( 3091 3082 )  100.n
R_D52311LOADxxQSG9 ( 3091 0 ) COMPLEX( 168.96,-126.72)
R_D52312xxQSG9 ( 3090 3082 )  100.n
R_D52312LOADxxQSG9 ( 3090 0 ) COMPLEX( 86.7843,-60.576)
R_D52313xxQSG9 ( 3089 3082 )  100.n
R_D52313LOADxxQSG9 ( 3089 0 ) COMPLEX( 6.078,-3.2805)
R_D52314xxQSG9 ( 3088 3082 )  100.n
R_D52314LOADxxQSG9 ( 3088 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG9 ( 3087 3082 )  100.n
R_D52315LOADxxQSG9 ( 3087 0 ) COMPLEX( 390., 0.)
R_D52316xxQSG9 ( 3086 3082 )  100.n
R_D52316LOADxxQSG9 ( 3086 0 ) COMPLEX( 10.7391,-6.372)
R_D52317xxQSG9 ( 3085 3082 )  100.n
R_D52317LOADxxQSG9 ( 3085 0 ) COMPLEX( 10.7391,-6.372)
R_D52310xxQSG9 ( 3084 3082 )  100.n
R_D52310LOADxxQSG9 ( 3084 0 ) COMPLEX( 168.96,-126.72)
R_D52309LOADxxQSG9 ( 0 3083 ) COMPLEX( 390., 0.)
R_D52309xxQSG9 ( 3083 3082 )  100.n
R_D52307LOADxxQSG9 ( 3081 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG9 ( 3081 3082 )  100.n
R_D52201xxQSG9 ( 3067 3080 )  100.n
R_D52201LOADxxQSG9 ( 0 3080 ) COMPLEX( 1.9074,-1.182)
R_D52202xxQSG9 ( 3079 3067 )  100.n
R_D52202LOADxxQSG9 ( 0 3079 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG9 ( 3078 3067 )  100.n
R_D52203LOADxxQSG9 ( 0 3078 ) COMPLEX( 390., 0.)
R_D52204xxQSG9 ( 3077 3067 )  100.n
R_D52204LOADxxQSG9 ( 0 3077 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG9 ( 3076 3067 )  100.n
R_D52205LOADxxQSG9 ( 0 3076 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG9 ( 3075 3067 )  100.n
R_D52206LOADxxQSG9 ( 3065 3075 )  100.n
R_D52208LOADxxQSG9 ( 0 3074 ) COMPLEX( 10.7391,-6.372)
R_D52208xxQSG9 ( 3074 3067 )  100.n
R_D52211xxQSG9 ( 3073 3067 )  100.n
R_D52211LOADxxQSG9 ( 3073 0 ) COMPLEX( 418.2288,-214.2651)
R_D52212xxQSG9 ( 3072 3067 )  100.n
R_D52212LOADxxQSG9 ( 3072 0 ) COMPLEX( 8.1777,-4.4139)
R_D52213xxQSG9 ( 3071 3067 )  100.n
R_D52213LOADxxQSG9 ( 3071 0 ) COMPLEX( 390., 0.)
R_D52214xxQSG9 ( 3070 3067 )  100.n
R_D52214LOADxxQSG9 ( 3070 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG9 ( 3069 3067 )  100.n
R_D52210LOADxxQSG9 ( 3069 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG9 ( 0 3068 ) COMPLEX( 390., 0.)
R_D52209xxQSG9 ( 3068 3067 )  100.n
R_D52207LOADxxQSG9 ( 3066 0 ) COMPLEX( 235.5726,-188.9955)
R_D52207xxQSG9 ( 3066 3067 )  100.n
R_D52114xxQSG9 ( 3063 3064 )  100.n
R_D52114LOADxxQSG9 ( 3063 0 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG10 
R_D52101xxQSG10 ( 3116 3174 )  100.n
R_D52101LOADxxQSG10 ( 0 3174 ) COMPLEX( 390., 0.)
R_D52102xxQSG10 ( 3173 3116 )  100.n
R_D52102LOADxxQSG10 ( 0 3173 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG10 ( 3172 3116 )  100.n
R_D52103LOADxxQSG10 ( 0 3172 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG10 ( 3171 3116 )  100.n
R_D52104LOADxxQSG10 ( 0 3171 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG10 ( 3170 3116 )  100.n
R_D52105LOADxxQSG10 ( 0 3170 ) COMPLEX( 390., 0.)
R_D52107xxQSG10 ( 3169 3116 )  100.n
R_D52107LOADxxQSG10 ( 0 3169 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSG10 ( 0 3168 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG10 ( 3168 3116 )  100.n
R_D52112xxQSG10 ( 3167 3116 )  100.n
R_D52112LOADxxQSG10 ( 3167 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG10 ( 3166 3116 )  100.n
R_D52113LOADxxQSG10 ( 3166 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG10 ( 3165 3116 )  100.n
R_D52114LOADxxQSG10 ( 3165 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG10 ( 3164 3116 )  100.n
R_D52115LOADxxQSG10 ( 3164 0 ) COMPLEX( 3.9963,-2.265)
R_D52116xxQSG10 ( 3163 3116 )  100.n
R_D52116LOADxxQSG10 ( 3163 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG10 ( 0 0 )  1.E+12
R_D52111xxQSG10 ( 3161 3116 )  100.n
R_D52111LOADxxQSG10 ( 3161 0 ) COMPLEX( 8.1777,-4.4139)
R_D52109LOADxxQSG10 ( 0 3160 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG10 ( 3160 3116 )  100.n
R_D52106LOADxxQSG10 ( 3158 3159 )  100.n
R_D52106xxQSG10 ( 3159 3116 )  100.n
R_D52L2xxQSG10 ( 3118 3143 )  100.n
R_D52E2xxQSG10 ( 492 3143 )  100.n
R_D52E1xxQSG10 ( 476 3116 )  100.n
R_D52201xxQSG10 ( 3143 3156 )  100.n
R_D52201LOADxxQSG10 ( 0 3156 ) COMPLEX( 42.4488,-29.6295)
R_D52202xxQSG10 ( 3155 3143 )  100.n
R_D52202LOADxxQSG10 ( 0 3155 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG10 ( 3154 3143 )  100.n
R_D52203LOADxxQSG10 ( 0 3154 ) COMPLEX( 390., 0.)
R_D52204xxQSG10 ( 3153 3143 )  100.n
R_D52204LOADxxQSG10 ( 0 3153 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG10 ( 3152 3143 )  100.n
R_D52205LOADxxQSG10 ( 0 3152 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG10 ( 3151 3143 )  100.n
R_D52206LOADxxQSG10 ( 3141 3151 )  100.n
R_D52208LOADxxQSG10 ( 0 3150 ) COMPLEX( 418.2288,-214.2651)
R_D52208xxQSG10 ( 3150 3143 )  100.n
R_D52211xxQSG10 ( 3149 3143 )  100.n
R_D52211LOADxxQSG10 ( 3149 0 ) COMPLEX( 418.2288,-214.2651)
R_D52212xxQSG10 ( 3148 3143 )  100.n
R_D52212LOADxxQSG10 ( 3148 0 ) COMPLEX( 8.1777,-4.4139)
R_D52213xxQSG10 ( 3147 3143 )  100.n
R_D52213LOADxxQSG10 ( 3147 0 ) COMPLEX( 390., 0.)
R_D52214xxQSG10 ( 3146 3143 )  100.n
R_D52214LOADxxQSG10 ( 3146 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG10 ( 3145 3143 )  100.n
R_D52210LOADxxQSG10 ( 3145 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG10 ( 0 3144 ) COMPLEX( 390., 0.)
R_D52209xxQSG10 ( 3144 3143 )  100.n
R_D52207LOADxxQSG10 ( 3142 0 ) COMPLEX( 235.5726,-188.9955)
R_D52207xxQSG10 ( 3142 3143 )  100.n
R_D52301xxQSG10 ( 3118 3140 )  100.n
R_D52301LOADxxQSG10 ( 0 3140 ) COMPLEX( 1.9074,-1.182)
R_D52302xxQSG10 ( 3139 3118 )  100.n
R_D52302LOADxxQSG10 ( 0 3139 ) COMPLEX( 1.7298,-0.9336)
R_D52303xxQSG10 ( 3138 3118 )  100.n
R_D52303LOADxxQSG10 ( 0 3138 ) COMPLEX( 390., 0.)
R_D52304xxQSG10 ( 3137 3118 )  100.n
R_D52304LOADxxQSG10 ( 0 3137 ) COMPLEX( 390., 0.)
R_D52305xxQSG10 ( 3136 3118 )  100.n
R_D52305LOADxxQSG10 ( 0 3136 ) COMPLEX( 390., 0.)
R_D52306xxQSG10 ( 3135 3118 )  100.n
R_D52306LOADxxQSG10 ( 0 3135 ) COMPLEX( 176.6793,-141.7467)
R_D52308LOADxxQSG10 ( 0 3134 ) COMPLEX( 2.4495,-0.8052)
R_D52308xxQSG10 ( 3134 3118 )  100.n
R_D52311xxQSG10 ( 3133 3118 )  100.n
R_D52311LOADxxQSG10 ( 3133 0 ) COMPLEX( 168.96,-126.72)
R_D52312xxQSG10 ( 3132 3118 )  100.n
R_D52312LOADxxQSG10 ( 3132 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG10 ( 3131 3118 )  100.n
R_D52313LOADxxQSG10 ( 3131 0 ) COMPLEX( 86.7843,-60.576)
R_D52314xxQSG10 ( 3130 3118 )  100.n
R_D52314LOADxxQSG10 ( 3130 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG10 ( 3129 3118 )  100.n
R_D52315LOADxxQSG10 ( 3129 0 ) COMPLEX( 6.078,-3.2805)
R_D52316xxQSG10 ( 3128 3118 )  100.n
R_D52316LOADxxQSG10 ( 3128 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG10 ( 3127 3118 )  100.n
R_D52317LOADxxQSG10 ( 3127 0 ) COMPLEX( 10.7391,-6.372)
R_D52310xxQSG10 ( 3126 3118 )  100.n
R_D52310LOADxxQSG10 ( 3126 0 ) COMPLEX( 390., 0.)
R_D52318xxQSG10 ( 3125 3118 )  100.n
R_D52318LOADxxQSG10 ( 3125 0 ) COMPLEX( 10.7391,-6.372)
R_D52319xxQSG10 ( 3124 3118 )  100.n
R_D52319LOADxxQSG10 ( 3124 0 ) COMPLEX( 355.0272,-247.8105)
R_D52309LOADxxQSG10 ( 0 3123 ) COMPLEX( 390., 0.)
R_D52309xxQSG10 ( 3123 3118 )  100.n
R_D52307LOADxxQSG10 ( 3122 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG10 ( 3122 3118 )  100.n
R_D52320xxQSG10 ( 3118 3121 )  100.n
R_D52320LOADxxQSG10 ( 0 3121 ) COMPLEX( 4.773,-2.832)
R_D52321xxQSG10 ( 3120 3118 )  100.n
R_D52321LOADxxQSG10 ( 0 3120 ) COMPLEX( 4.773,-2.832)
R_D52323xxQSG10 ( 3119 3118 )  100.n
R_D52323LOADxxQSG10 ( 3119 0 ) COMPLEX( 2.322,-1.3779)
R_D52322xxQSG10 ( 3117 3118 )  100.n
R_D52322LOADxxQSG10 ( 3117 0 ) COMPLEX( 21.6276,-14.5338)
R_D52110LOADxxQSG10 ( 0 3115 ) COMPLEX( 418.2288,-214.2651)
R_D52110xxQSG10 ( 3115 3116 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG11 
R_D52101xxQSG11 ( 3176 3234 )  100.n
R_D52101LOADxxQSG11 ( 0 3234 ) COMPLEX( 102.99,-74.5635)
R_D52102xxQSG11 ( 3233 3176 )  100.n
R_D52102LOADxxQSG11 ( 0 3233 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG11 ( 3232 3176 )  100.n
R_D52103LOADxxQSG11 ( 0 3232 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG11 ( 3231 3176 )  100.n
R_D52104LOADxxQSG11 ( 0 3231 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG11 ( 3230 3176 )  100.n
R_D52105LOADxxQSG11 ( 0 3230 ) COMPLEX( 390., 0.)
R_D52106xxQSG11 ( 3229 3176 )  100.n
R_D52106LOADxxQSG11 ( 0 3229 ) COMPLEX( 4.773,-2.832)
R_D52108LOADxxQSG11 ( 0 3228 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG11 ( 3228 3176 )  100.n
R_D52112xxQSG11 ( 3227 3176 )  100.n
R_D52112LOADxxQSG11 ( 3227 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG11 ( 3226 3176 )  100.n
R_D52113LOADxxQSG11 ( 3226 0 ) COMPLEX( 3.9963,-2.265)
R_D52114xxQSG11 ( 3225 3176 )  100.n
R_D52114LOADxxQSG11 ( 3225 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG11 ( 3224 3176 )  100.n
R_D52115LOADxxQSG11 ( 3224 0 ) COMPLEX( 3.9963,-2.265)
R_D52116xxQSG11 ( 3223 3176 )  100.n
R_D52116LOADxxQSG11 ( 3223 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG11 ( 0 0 )  1.E+12
R_D52111xxQSG11 ( 3221 3176 )  100.n
R_D52111LOADxxQSG11 ( 3221 0 ) COMPLEX( 8.1777,-4.4139)
R_D52109LOADxxQSG11 ( 0 3220 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG11 ( 3220 3176 )  100.n
R_D52107LOADxxQSG11 ( 0 0 )  1.E+12
R_D52107xxQSG11 ( 3219 3176 )  100.n
R_D52L2xxQSG11 ( 3178 3203 )  100.n
R_D52E2xxQSG11 ( 405 3203 )  100.n
R_D52E1xxQSG11 ( 534 3176 )  100.n
R_D52201xxQSG11 ( 3203 3216 )  100.n
R_D52201LOADxxQSG11 ( 0 3216 ) COMPLEX( 42.4488,-29.6295)
R_D52202xxQSG11 ( 3215 3203 )  100.n
R_D52202LOADxxQSG11 ( 0 3215 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG11 ( 3214 3203 )  100.n
R_D52203LOADxxQSG11 ( 0 3214 ) COMPLEX( 390., 0.)
R_D52204xxQSG11 ( 3213 3203 )  100.n
R_D52204LOADxxQSG11 ( 0 3213 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG11 ( 3212 3203 )  100.n
R_D52205LOADxxQSG11 ( 0 3212 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG11 ( 3211 3203 )  100.n
R_D52206LOADxxQSG11 ( 0 0 )  1.E+12
R_D52208LOADxxQSG11 ( 0 3210 ) COMPLEX( 4.773,-2.832)
R_D52208xxQSG11 ( 3210 3203 )  100.n
R_D52211xxQSG11 ( 3209 3203 )  100.n
R_D52211LOADxxQSG11 ( 3209 0 ) COMPLEX( 418.2288,-214.2651)
R_D52212xxQSG11 ( 3208 3203 )  100.n
R_D52212LOADxxQSG11 ( 3208 0 ) COMPLEX( 8.1777,-4.4139)
R_D52213xxQSG11 ( 3207 3203 )  100.n
R_D52213LOADxxQSG11 ( 3207 0 ) COMPLEX( 13.9875,-8.6688)
R_D52214xxQSG11 ( 3206 3203 )  100.n
R_D52214LOADxxQSG11 ( 3206 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG11 ( 3205 3203 )  100.n
R_D52210LOADxxQSG11 ( 3205 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG11 ( 0 3204 ) COMPLEX( 3.9963,-2.265)
R_D52209xxQSG11 ( 3204 3203 )  100.n
R_D52207LOADxxQSG11 ( 3202 0 ) COMPLEX( 235.5726,-188.9955)
R_D52207xxQSG11 ( 3202 3203 )  100.n
R_D52301xxQSG11 ( 3178 3200 )  100.n
R_D52301LOADxxQSG11 ( 0 3200 ) COMPLEX( 1.9074,-1.182)
R_D52302xxQSG11 ( 3199 3178 )  100.n
R_D52302LOADxxQSG11 ( 0 3199 ) COMPLEX( 1.2714,-0.6159)
R_D52303xxQSG11 ( 3198 3178 )  100.n
R_D52303LOADxxQSG11 ( 0 3198 ) COMPLEX( 390., 0.)
R_D52304xxQSG11 ( 3197 3178 )  100.n
R_D52304LOADxxQSG11 ( 0 3197 ) COMPLEX( 176.6793,-141.7467)
R_D52305xxQSG11 ( 3196 3178 )  100.n
R_D52305LOADxxQSG11 ( 0 3196 ) COMPLEX( 168.96,-126.72)
R_D52306xxQSG11 ( 3195 3178 )  100.n
R_D52306LOADxxQSG11 ( 0 3195 ) COMPLEX( 390., 0.)
R_D52308LOADxxQSG11 ( 0 3194 ) COMPLEX( 2.4495,-0.8052)
R_D52308xxQSG11 ( 3194 3178 )  100.n
R_D52311xxQSG11 ( 3193 3178 )  100.n
R_D52311LOADxxQSG11 ( 3193 0 ) COMPLEX( 168.96,-126.72)
R_D52312xxQSG11 ( 3192 3178 )  100.n
R_D52312LOADxxQSG11 ( 3192 0 ) COMPLEX( 168.96,-126.72)
R_D52313xxQSG11 ( 3191 3178 )  100.n
R_D52313LOADxxQSG11 ( 3191 0 ) COMPLEX( 86.7843,-60.576)
R_D52314xxQSG11 ( 3190 3178 )  100.n
R_D52314LOADxxQSG11 ( 3190 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG11 ( 3189 3178 )  100.n
R_D52315LOADxxQSG11 ( 3189 0 ) COMPLEX( 6.078,-3.2805)
R_D52316xxQSG11 ( 3188 3178 )  100.n
R_D52316LOADxxQSG11 ( 3188 0 ) COMPLEX( 390., 0.)
R_D52317xxQSG11 ( 3187 3178 )  100.n
R_D52317LOADxxQSG11 ( 3187 0 ) COMPLEX( 10.7391,-6.372)
R_D52310xxQSG11 ( 3186 3178 )  100.n
R_D52310LOADxxQSG11 ( 3186 0 ) COMPLEX( 6.078,-3.2805)
R_D52318xxQSG11 ( 3185 3178 )  100.n
R_D52318LOADxxQSG11 ( 3185 0 ) COMPLEX( 10.7391,-6.372)
R_D52319xxQSG11 ( 3184 3178 )  100.n
R_D52319LOADxxQSG11 ( 3184 0 ) COMPLEX( 6.078,-3.2805)
R_D52309LOADxxQSG11 ( 0 3183 ) COMPLEX( 390., 0.)
R_D52309xxQSG11 ( 3183 3178 )  100.n
R_D52307LOADxxQSG11 ( 3182 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG11 ( 3182 3178 )  100.n
R_D52320xxQSG11 ( 3178 3181 )  100.n
R_D52320LOADxxQSG11 ( 0 3181 ) COMPLEX( 4.2531,-2.5236)
R_D52321xxQSG11 ( 3180 3178 )  100.n
R_D52321LOADxxQSG11 ( 0 3180 ) COMPLEX( 390., 0.)
R_D52323xxQSG11 ( 3179 3178 )  100.n
R_D52323LOADxxQSG11 ( 3179 0 ) COMPLEX( 2.4495,-0.8052)
R_D52322xxQSG11 ( 3177 3178 )  100.n
R_D52322LOADxxQSG11 ( 3177 0 ) COMPLEX( 21.6276,-14.5338)
R_D52110LOADxxQSG11 ( 0 3175 ) COMPLEX( 418.2288,-214.2651)
R_D52110xxQSG11 ( 3175 3176 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG12 
R_D52101xxQSG12 ( 3236 3289 )  100.n
R_D52101LOADxxQSG12 ( 0 3289 ) COMPLEX( 390., 0.)
R_D52102xxQSG12 ( 3288 3236 )  100.n
R_D52102LOADxxQSG12 ( 0 3288 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG12 ( 3287 3236 )  100.n
R_D52103LOADxxQSG12 ( 0 3287 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG12 ( 3286 3236 )  100.n
R_D52104LOADxxQSG12 ( 0 3286 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG12 ( 3285 3236 )  100.n
R_D52105LOADxxQSG12 ( 0 3285 ) COMPLEX( 390., 0.)
R_D52106xxQSG12 ( 3284 3236 )  100.n
R_D52106LOADxxQSG12 ( 3273 3284 )  100.n
R_D52108LOADxxQSG12 ( 0 3283 ) COMPLEX( 3.9963,-2.265)
R_D52108xxQSG12 ( 3283 3236 )  100.n
R_D52112xxQSG12 ( 3282 3236 )  100.n
R_D52112LOADxxQSG12 ( 3282 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG12 ( 3281 3236 )  100.n
R_D52113LOADxxQSG12 ( 3281 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG12 ( 3280 3236 )  100.n
R_D52114LOADxxQSG12 ( 3280 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG12 ( 3279 3236 )  100.n
R_D52115LOADxxQSG12 ( 3279 0 ) COMPLEX( 3.9963,-2.265)
R_D52116xxQSG12 ( 3278 3236 )  100.n
R_D52116LOADxxQSG12 ( 3278 0 ) COMPLEX( 3.9963,-2.265)
R_D52L1xxQSG12 ( 0 0 )  1.E+12
R_D52111xxQSG12 ( 3276 3236 )  100.n
R_D52111LOADxxQSG12 ( 3276 0 ) COMPLEX( 8.1777,-4.4139)
R_D52109LOADxxQSG12 ( 0 3275 ) COMPLEX( 3.9963,-2.265)
R_D52109xxQSG12 ( 3275 3236 )  100.n
R_D52107LOADxxQSG12 ( 3274 0 ) COMPLEX( 390., 0.)
R_D52107xxQSG12 ( 3274 3236 )  100.n
R_D52L2xxQSG12 ( 3254 3239 )  100.n
R_D52E2xxQSG12 ( 541 3239 )  100.n
R_D52E1xxQSG12 ( 409 3236 )  100.n
R_D52301xxQSG12 ( 3254 3271 )  100.n
R_D52301LOADxxQSG12 ( 0 3271 ) COMPLEX( 1.9074,-1.182)
R_D52302xxQSG12 ( 3270 3254 )  100.n
R_D52302LOADxxQSG12 ( 0 3270 ) COMPLEX( 390., 0.)
R_D52303xxQSG12 ( 3269 3254 )  100.n
R_D52303LOADxxQSG12 ( 0 3269 ) COMPLEX( 390., 0.)
R_D52304xxQSG12 ( 3268 3254 )  100.n
R_D52304LOADxxQSG12 ( 0 3268 ) COMPLEX( 390., 0.)
R_D52305xxQSG12 ( 3267 3254 )  100.n
R_D52305LOADxxQSG12 ( 0 3267 ) COMPLEX( 390., 0.)
R_D52306xxQSG12 ( 3266 3254 )  100.n
R_D52306LOADxxQSG12 ( 0 3266 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG12 ( 0 3265 ) COMPLEX( 390., 0.)
R_D52308xxQSG12 ( 3265 3254 )  100.n
R_D52311xxQSG12 ( 3264 3254 )  100.n
R_D52311LOADxxQSG12 ( 3264 0 ) COMPLEX( 168.96,-126.72)
R_D52312xxQSG12 ( 3263 3254 )  100.n
R_D52312LOADxxQSG12 ( 3263 0 ) COMPLEX( 86.7843,-60.576)
R_D52313xxQSG12 ( 3262 3254 )  100.n
R_D52313LOADxxQSG12 ( 3262 0 ) COMPLEX( 6.078,-3.2805)
R_D52314xxQSG12 ( 3261 3254 )  100.n
R_D52314LOADxxQSG12 ( 3261 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG12 ( 3260 3254 )  100.n
R_D52315LOADxxQSG12 ( 3260 0 ) COMPLEX( 390., 0.)
R_D52316xxQSG12 ( 3259 3254 )  100.n
R_D52316LOADxxQSG12 ( 3259 0 ) COMPLEX( 10.7391,-6.372)
R_D52317xxQSG12 ( 3258 3254 )  100.n
R_D52317LOADxxQSG12 ( 3258 0 ) COMPLEX( 10.7391,-6.372)
R_D52310xxQSG12 ( 3257 3254 )  100.n
R_D52310LOADxxQSG12 ( 3257 0 ) COMPLEX( 168.96,-126.72)
R_D52318xxQSG12 ( 3256 3254 )  100.n
R_D52318LOADxxQSG12 ( 3256 0 ) COMPLEX( 176.6793,-141.7467)
R_D52309LOADxxQSG12 ( 0 3255 ) COMPLEX( 390., 0.)
R_D52309xxQSG12 ( 3255 3254 )  100.n
R_D52307LOADxxQSG12 ( 3253 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG12 ( 3253 3254 )  100.n
R_D52201xxQSG12 ( 3239 3252 )  100.n
R_D52201LOADxxQSG12 ( 0 3252 ) COMPLEX( 42.4488,-29.6295)
R_D52202xxQSG12 ( 3251 3239 )  100.n
R_D52202LOADxxQSG12 ( 0 3251 ) COMPLEX( 86.7843,-60.576)
R_D52203xxQSG12 ( 3250 3239 )  100.n
R_D52203LOADxxQSG12 ( 0 3250 ) COMPLEX( 390., 0.)
R_D52204xxQSG12 ( 3249 3239 )  100.n
R_D52204LOADxxQSG12 ( 0 3249 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG12 ( 3248 3239 )  100.n
R_D52205LOADxxQSG12 ( 0 3248 ) COMPLEX( 3.9963,-2.265)
R_D52206xxQSG12 ( 3247 3239 )  100.n
R_D52206LOADxxQSG12 ( 3237 3247 )  100.n
R_D52208LOADxxQSG12 ( 0 3246 ) COMPLEX( 390., 0.)
R_D52208xxQSG12 ( 3246 3239 )  100.n
R_D52211xxQSG12 ( 3245 3239 )  100.n
R_D52211LOADxxQSG12 ( 3245 0 ) COMPLEX( 418.2288,-214.2651)
R_D52212xxQSG12 ( 3244 3239 )  100.n
R_D52212LOADxxQSG12 ( 3244 0 ) COMPLEX( 8.1777,-4.4139)
R_D52213xxQSG12 ( 3243 3239 )  100.n
R_D52213LOADxxQSG12 ( 3243 0 ) COMPLEX( 390., 0.)
R_D52214xxQSG12 ( 3242 3239 )  100.n
R_D52214LOADxxQSG12 ( 3242 0 ) COMPLEX( 3.9963,-2.265)
R_D52210xxQSG12 ( 3241 3239 )  100.n
R_D52210LOADxxQSG12 ( 3241 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG12 ( 0 3240 ) COMPLEX( 390., 0.)
R_D52209xxQSG12 ( 3240 3239 )  100.n
R_D52207LOADxxQSG12 ( 3238 0 ) COMPLEX( 235.5726,-188.9955)
R_D52207xxQSG12 ( 3238 3239 )  100.n
R_D52110LOADxxQSG12 ( 0 3235 ) COMPLEX( 418.2288,-214.2651)
R_D52110xxQSG12 ( 3235 3236 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSG13 
R_D52101xxQSG13 ( 3291 3341 )  100.n
R_D52101LOADxxQSG13 ( 0 3341 ) COMPLEX( 53.3484,-35.8503)
R_D52102xxQSG13 ( 3340 3291 )  100.n
R_D52102LOADxxQSG13 ( 0 3340 ) COMPLEX( 86.7843,-60.576)
R_D52103xxQSG13 ( 3339 3291 )  100.n
R_D52103LOADxxQSG13 ( 0 3339 ) COMPLEX( 3.9963,-2.265)
R_D52104xxQSG13 ( 3338 3291 )  100.n
R_D52104LOADxxQSG13 ( 0 3338 ) COMPLEX( 3.9963,-2.265)
R_D52105xxQSG13 ( 3337 3291 )  100.n
R_D52105LOADxxQSG13 ( 0 3337 ) COMPLEX( 390., 0.)
R_D52106xxQSG13 ( 3336 3291 )  100.n
R_D52106LOADxxQSG13 ( 0 3336 ) COMPLEX( 102.99,-74.5635)
R_D52108LOADxxQSG13 ( 0 3335 ) COMPLEX( 390., 0.)
R_D52108xxQSG13 ( 3335 3291 )  100.n
R_D52112xxQSG13 ( 3334 3291 )  100.n
R_D52112LOADxxQSG13 ( 3334 0 ) COMPLEX( 390., 0.)
R_D52113xxQSG13 ( 3333 3291 )  100.n
R_D52113LOADxxQSG13 ( 3333 0 ) COMPLEX( 390., 0.)
R_D52114xxQSG13 ( 3332 3291 )  100.n
R_D52114LOADxxQSG13 ( 3332 0 ) COMPLEX( 390., 0.)
R_D52115xxQSG13 ( 3331 3291 )  100.n
R_D52115LOADxxQSG13 ( 3331 0 ) COMPLEX( 2.322,-1.3779)
R_D52L1xxQSG13 ( 0 0 )  1.E+12
R_D52111xxQSG13 ( 3329 3291 )  100.n
R_D52111LOADxxQSG13 ( 3329 0 ) COMPLEX( 8.1777,-4.4139)
R_D52109LOADxxQSG13 ( 0 3328 ) COMPLEX( 390., 0.)
R_D52109xxQSG13 ( 3328 3291 )  100.n
R_D52107LOADxxQSG13 ( 3327 0 ) COMPLEX( 390., 0.)
R_D52107xxQSG13 ( 3327 3291 )  100.n
R_D52L2xxQSG13 ( 3308 3293 )  100.n
R_D52E2xxQSG13 ( 397 3293 )  100.n
R_D52E1xxQSG13 ( 414 3291 )  100.n
R_D52301xxQSG13 ( 3308 3325 )  100.n
R_D52301LOADxxQSG13 ( 0 3325 ) COMPLEX( 390., 0.)
R_D52302xxQSG13 ( 3324 3308 )  100.n
R_D52302LOADxxQSG13 ( 0 3324 ) COMPLEX( 390., 0.)
R_D52303xxQSG13 ( 3323 3308 )  100.n
R_D52303LOADxxQSG13 ( 0 3323 ) COMPLEX( 235.5726,-188.9955)
R_D52304xxQSG13 ( 3322 3308 )  100.n
R_D52304LOADxxQSG13 ( 0 3322 ) COMPLEX( 30.976, 0.)
R_D52305xxQSG13 ( 3321 3308 )  100.n
R_D52305LOADxxQSG13 ( 0 3321 ) COMPLEX( 390., 0.)
R_D52306xxQSG13 ( 3320 3308 )  100.n
R_D52306LOADxxQSG13 ( 0 3320 ) COMPLEX( 2.4495,-0.8052)
R_D52308LOADxxQSG13 ( 0 3319 ) COMPLEX( 10.9203,-3.5892)
R_D52308xxQSG13 ( 3319 3308 )  100.n
R_D52311xxQSG13 ( 3318 3308 )  100.n
R_D52311LOADxxQSG13 ( 3318 0 ) COMPLEX( 168.96,-126.72)
R_D52312xxQSG13 ( 3317 3308 )  100.n
R_D52312LOADxxQSG13 ( 3317 0 ) COMPLEX( 390., 0.)
R_D52313xxQSG13 ( 3316 3308 )  100.n
R_D52313LOADxxQSG13 ( 3316 0 ) COMPLEX( 6.078,-3.2805)
R_D52314xxQSG13 ( 3315 3308 )  100.n
R_D52314LOADxxQSG13 ( 3315 0 ) COMPLEX( 6.078,-3.2805)
R_D52315xxQSG13 ( 3314 3308 )  100.n
R_D52315LOADxxQSG13 ( 3314 0 ) COMPLEX( 390., 0.)
R_D52316xxQSG13 ( 3313 3308 )  100.n
R_D52316LOADxxQSG13 ( 3313 0 ) COMPLEX( 10.7391,-6.372)
R_D52317xxQSG13 ( 3312 3308 )  100.n
R_D52317LOADxxQSG13 ( 3312 0 ) COMPLEX( 10.7391,-6.372)
R_D52310xxQSG13 ( 3311 3308 )  100.n
R_D52310LOADxxQSG13 ( 3311 0 ) COMPLEX( 168.96,-126.72)
R_D52318xxQSG13 ( 3310 3308 )  100.n
R_D52318LOADxxQSG13 ( 3310 0 ) COMPLEX( 176.6793,-141.7467)
R_D52309LOADxxQSG13 ( 0 3309 ) COMPLEX( 390., 0.)
R_D52309xxQSG13 ( 3309 3308 )  100.n
R_D52307LOADxxQSG13 ( 3307 0 ) COMPLEX( 2.4495,-0.8052)
R_D52307xxQSG13 ( 3307 3308 )  100.n
R_D52201xxQSG13 ( 3293 3306 )  100.n
R_D52201LOADxxQSG13 ( 0 3306 ) COMPLEX( 390., 0.)
R_D52202xxQSG13 ( 3305 3293 )  100.n
R_D52202LOADxxQSG13 ( 0 3305 ) COMPLEX( 390., 0.)
R_D52203xxQSG13 ( 3304 3293 )  100.n
R_D52203LOADxxQSG13 ( 0 3304 ) COMPLEX( 390., 0.)
R_D52204xxQSG13 ( 3303 3293 )  100.n
R_D52204LOADxxQSG13 ( 0 3303 ) COMPLEX( 3.9963,-2.265)
R_D52205xxQSG13 ( 3302 3293 )  100.n
R_D52205LOADxxQSG13 ( 0 3302 ) COMPLEX( 390., 0.)
R_D52206xxQSG13 ( 3301 3293 )  100.n
R_D52206LOADxxQSG13 ( 0 3301 ) COMPLEX( 390., 0.)
R_D52208LOADxxQSG13 ( 0 3300 ) COMPLEX( 390., 0.)
R_D52208xxQSG13 ( 3300 3293 )  100.n
R_D52211xxQSG13 ( 3299 3293 )  100.n
R_D52211LOADxxQSG13 ( 3299 0 ) COMPLEX( 418.2288,-214.2651)
R_D52212xxQSG13 ( 3298 3293 )  100.n
R_D52212LOADxxQSG13 ( 3298 0 ) COMPLEX( 8.1777,-4.4139)
R_D52213xxQSG13 ( 3297 3293 )  100.n
R_D52213LOADxxQSG13 ( 3297 0 ) COMPLEX( 390., 0.)
R_D52214xxQSG13 ( 3296 3293 )  100.n
R_D52214LOADxxQSG13 ( 3296 0 ) COMPLEX( 2.322,-1.3779)
R_D52210xxQSG13 ( 3295 3293 )  100.n
R_D52210LOADxxQSG13 ( 3295 0 ) COMPLEX( 390., 0.)
R_D52209LOADxxQSG13 ( 0 3294 ) COMPLEX( 390., 0.)
R_D52209xxQSG13 ( 3294 3293 )  100.n
R_D52207LOADxxQSG13 ( 3292 0 ) COMPLEX( 390., 0.)
R_D52207xxQSG13 ( 3292 3293 )  100.n
R_D52110LOADxxQSG13 ( 0 3290 ) COMPLEX( 418.2288,-214.2651)
R_D52110xxQSG13 ( 3290 3291 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE8 
R_D52E1xxQSSE8 ( 604 3347 )  100.n
R_D52E2xxQSSE8 ( 485 3351 )  100.n
R_D52306xxQSSE8 ( 3360 3343 )  100.n
R_D52306LOADxxQSSE8 ( 0 3360 ) COMPLEX( 390., 0.)
R_D52104xxQSSE8 ( 3359 3347 )  100.n
R_D52104LOADxxQSSE8 ( 0 3359 ) COMPLEX( 390., 0.)
R_D52305xxQSSE8 ( 3358 3343 )  100.n
R_D52305LOADxxQSSE8 ( 0 3358 ) COMPLEX( 11.6484,-3.8286)
R_D52304xxQSSE8 ( 3357 3343 )  100.n
R_D52304LOADxxQSSE8 ( 0 3357 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE8 ( 3356 3343 )  100.n
R_D52303LOADxxQSSE8 ( 0 3356 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE8 ( 3355 3343 )  100.n
R_D52302LOADxxQSSE8 ( 0 3355 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE8 ( 3354 3343 )  100.n
R_D52301LOADxxQSSE8 ( 0 3354 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE8 ( 3353 3351 )  100.n
R_D52203LOADxxQSSE8 ( 0 3353 ) COMPLEX( 390., 0.)
R_D52202xxQSSE8 ( 3352 3351 )  100.n
R_D52202LOADxxQSSE8 ( 0 3352 ) COMPLEX( 390., 0.)
R_D52201xxQSSE8 ( 3350 3351 )  100.n
R_D52201LOADxxQSSE8 ( 0 3350 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE8 ( 3349 3347 )  100.n
R_D52103LOADxxQSSE8 ( 0 3349 ) COMPLEX( 390., 0.)
R_D52102xxQSSE8 ( 3348 3347 )  100.n
R_D52102LOADxxQSSE8 ( 0 3348 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE8 ( 3346 3347 )  100.n
R_D52101LOADxxQSSE8 ( 0 3346 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE8 ( 0 0 )  1.E+12
R_D52L2xxQSSE8 ( 3343 3351 )  100.n
R_D52309xxQSSE8 ( 3345 3343 )  100.n
R_D52309LOADxxQSSE8 ( 0 3345 ) COMPLEX( 390., 0.)
R_D52308xxQSSE8 ( 3344 3343 )  100.n
R_D52308LOADxxQSSE8 ( 0 3344 ) COMPLEX( 390., 0.)
R_D52307xxQSSE8 ( 3342 3343 )  100.n
R_D52307LOADxxQSSE8 ( 0 3342 ) COMPLEX( 11.6484,-3.8286)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE9 
R_D52E1xxQSSE9 ( 488 3363 )  100.n
R_D52E2xxQSSE9 ( 612 3367 )  100.n
R_D52307xxQSSE9 ( 3376 3361 )  100.n
R_D52307LOADxxQSSE9 ( 0 3376 ) COMPLEX( 390., 0.)
R_D52306xxQSSE9 ( 3375 3361 )  100.n
R_D52306LOADxxQSSE9 ( 0 3375 ) COMPLEX( 390., 0.)
R_D52305xxQSSE9 ( 3374 3361 )  100.n
R_D52305LOADxxQSSE9 ( 0 3374 ) COMPLEX( 390., 0.)
R_D52304xxQSSE9 ( 3373 3361 )  100.n
R_D52304LOADxxQSSE9 ( 0 3373 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE9 ( 3372 3361 )  100.n
R_D52303LOADxxQSSE9 ( 0 3372 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE9 ( 3371 3361 )  100.n
R_D52302LOADxxQSSE9 ( 0 3371 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE9 ( 3370 3361 )  100.n
R_D52301LOADxxQSSE9 ( 0 3370 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE9 ( 3369 3367 )  100.n
R_D52203LOADxxQSSE9 ( 0 3369 ) COMPLEX( 390., 0.)
R_D52202xxQSSE9 ( 3368 3367 )  100.n
R_D52202LOADxxQSSE9 ( 0 3368 ) COMPLEX( 390., 0.)
R_D52201xxQSSE9 ( 3366 3367 )  100.n
R_D52201LOADxxQSSE9 ( 0 3366 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE9 ( 3365 3363 )  100.n
R_D52103LOADxxQSSE9 ( 0 3365 ) COMPLEX( 390., 0.)
R_D52102xxQSSE9 ( 3364 3363 )  100.n
R_D52102LOADxxQSSE9 ( 0 3364 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE9 ( 3362 3363 )  100.n
R_D52101LOADxxQSSE9 ( 0 3362 ) COMPLEX( 390., 0.)
R_D52L1xxQSSE9 ( 0 0 )  1.E+12
R_D52L2xxQSSE9 ( 3361 3367 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE10 
R_D52E1xxQSSE10 ( 477 3382 )  100.n
R_D52E2xxQSSE10 ( 496 3386 )  100.n
R_D52104xxQSSE10 ( 3394 3382 )  100.n
R_D52104LOADxxQSSE10 ( 0 3394 ) COMPLEX( 390., 0.)
R_D52305xxQSSE10 ( 3393 3378 )  100.n
R_D52305LOADxxQSSE10 ( 0 3393 ) COMPLEX( 11.6484,-3.8286)
R_D52304xxQSSE10 ( 3392 3378 )  100.n
R_D52304LOADxxQSSE10 ( 0 3392 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE10 ( 3391 3378 )  100.n
R_D52303LOADxxQSSE10 ( 0 3391 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE10 ( 3390 3378 )  100.n
R_D52302LOADxxQSSE10 ( 0 3390 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE10 ( 3389 3378 )  100.n
R_D52301LOADxxQSSE10 ( 0 3389 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE10 ( 3388 3386 )  100.n
R_D52203LOADxxQSSE10 ( 0 3388 ) COMPLEX( 390., 0.)
R_D52202xxQSSE10 ( 3387 3386 )  100.n
R_D52202LOADxxQSSE10 ( 0 3387 ) COMPLEX( 390., 0.)
R_D52201xxQSSE10 ( 3385 3386 )  100.n
R_D52201LOADxxQSSE10 ( 0 3385 ) COMPLEX( 30.976, 0.)
R_D52103xxQSSE10 ( 3384 3382 )  100.n
R_D52103LOADxxQSSE10 ( 0 3384 ) COMPLEX( 161.6139,-121.2105)
R_D52102xxQSSE10 ( 3383 3382 )  100.n
R_D52102LOADxxQSSE10 ( 0 3383 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE10 ( 3381 3382 )  100.n
R_D52101LOADxxQSSE10 ( 0 3381 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE10 ( 0 0 )  1.E+12
R_D52L2xxQSSE10 ( 3378 3386 )  100.n
R_D52306xxQSSE10 ( 3380 3378 )  100.n
R_D52306LOADxxQSSE10 ( 0 3380 ) COMPLEX( 390., 0.)
R_D52308xxQSSE10 ( 3379 3378 )  100.n
R_D52308LOADxxQSSE10 ( 0 3379 ) COMPLEX( 390., 0.)
R_D52307xxQSSE10 ( 3377 3378 )  100.n
R_D52307LOADxxQSSE10 ( 0 3377 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE11 
R_D52E1xxQSSE11 ( 535 3398 )  100.n
R_D52E2xxQSSE11 ( 395 3402 )  100.n
R_D52306xxQSSE11 ( 3410 3396 )  100.n
R_D52306LOADxxQSSE11 ( 0 3410 ) COMPLEX( 390., 0.)
R_D52305xxQSSE11 ( 3409 3396 )  100.n
R_D52305LOADxxQSSE11 ( 0 3409 ) COMPLEX( 11.6484,-3.8286)
R_D52304xxQSSE11 ( 3408 3396 )  100.n
R_D52304LOADxxQSSE11 ( 0 3408 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE11 ( 3407 3396 )  100.n
R_D52303LOADxxQSSE11 ( 0 3407 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE11 ( 3406 3396 )  100.n
R_D52302LOADxxQSSE11 ( 0 3406 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE11 ( 3405 3396 )  100.n
R_D52301LOADxxQSSE11 ( 0 3405 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE11 ( 3404 3402 )  100.n
R_D52203LOADxxQSSE11 ( 0 3404 ) COMPLEX( 390., 0.)
R_D52202xxQSSE11 ( 3403 3402 )  100.n
R_D52202LOADxxQSSE11 ( 0 3403 ) COMPLEX( 390., 0.)
R_D52201xxQSSE11 ( 3401 3402 )  100.n
R_D52201LOADxxQSSE11 ( 0 3401 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE11 ( 3400 3398 )  100.n
R_D52103LOADxxQSSE11 ( 0 3400 ) COMPLEX( 390., 0.)
R_D52102xxQSSE11 ( 3399 3398 )  100.n
R_D52102LOADxxQSSE11 ( 0 3399 ) COMPLEX( 390., 0.)
R_D52101xxQSSE11 ( 3397 3398 )  100.n
R_D52101LOADxxQSSE11 ( 0 3397 ) COMPLEX( 161.6139,-121.2105)
R_D52L1xxQSSE11 ( 0 0 )  1.E+12
R_D52L2xxQSSE11 ( 3396 3402 )  100.n
R_D52307xxQSSE11 ( 3395 3396 )  100.n
R_D52307LOADxxQSSE11 ( 0 3395 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE12 
R_D52E1xxQSSE12 ( 410 3412 )  100.n
R_D52E2xxQSSE12 ( 543 3419 )  100.n
R_D52306xxQSSE12 ( 3427 3414 )  100.n
R_D52306LOADxxQSSE12 ( 0 3427 ) COMPLEX( 390., 0.)
R_D52305xxQSSE12 ( 3426 3414 )  100.n
R_D52305LOADxxQSSE12 ( 0 3426 ) COMPLEX( 390., 0.)
R_D52304xxQSSE12 ( 3425 3414 )  100.n
R_D52304LOADxxQSSE12 ( 0 3425 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE12 ( 3424 3414 )  100.n
R_D52303LOADxxQSSE12 ( 0 3424 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE12 ( 3423 3414 )  100.n
R_D52302LOADxxQSSE12 ( 0 3423 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE12 ( 3422 3414 )  100.n
R_D52301LOADxxQSSE12 ( 0 3422 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE12 ( 3421 3419 )  100.n
R_D52203LOADxxQSSE12 ( 0 3421 ) COMPLEX( 390., 0.)
R_D52202xxQSSE12 ( 3420 3419 )  100.n
R_D52202LOADxxQSSE12 ( 0 3420 ) COMPLEX( 390., 0.)
R_D52201xxQSSE12 ( 3418 3419 )  100.n
R_D52201LOADxxQSSE12 ( 0 3418 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE12 ( 3417 3412 )  100.n
R_D52103LOADxxQSSE12 ( 0 3417 ) COMPLEX( 390., 0.)
R_D52102xxQSSE12 ( 3416 3412 )  100.n
R_D52102LOADxxQSSE12 ( 0 3416 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE12 ( 3415 3412 )  100.n
R_D52101LOADxxQSSE12 ( 0 3415 ) COMPLEX( 390., 0.)
R_D52L1xxQSSE12 ( 0 0 )  1.E+12
R_D52L2xxQSSE12 ( 3414 3419 )  100.n
R_D52307xxQSSE12 ( 3413 3414 )  100.n
R_D52307LOADxxQSSE12 ( 0 3413 ) COMPLEX( 390., 0.)
R_D52104xxQSSE12 ( 3411 3412 )  100.n
R_D52104LOADxxQSSE12 ( 0 3411 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSSE13 
R_D52E1xxQSSE13 ( 418 3431 )  100.n
R_D52E2xxQSSE13 ( 398 3437 )  100.n
R_D52306xxQSSE13 ( 3445 3429 )  100.n
R_D52306LOADxxQSSE13 ( 0 3445 ) COMPLEX( 11.6484,-3.8286)
R_D52305xxQSSE13 ( 3444 3429 )  100.n
R_D52305LOADxxQSSE13 ( 0 3444 ) COMPLEX( 390., 0.)
R_D52304xxQSSE13 ( 3443 3429 )  100.n
R_D52304LOADxxQSSE13 ( 0 3443 ) COMPLEX( 747.3483,-783.9678)
R_D52303xxQSSE13 ( 3442 3429 )  100.n
R_D52303LOADxxQSSE13 ( 0 3442 ) COMPLEX( 747.3483,-783.9678)
R_D52302xxQSSE13 ( 3441 3429 )  100.n
R_D52302LOADxxQSSE13 ( 0 3441 ) COMPLEX( 11.6484,-3.8286)
R_D52301xxQSSE13 ( 3440 3429 )  100.n
R_D52301LOADxxQSSE13 ( 0 3440 ) COMPLEX( 10.7391,-6.372)
R_D52203xxQSSE13 ( 3439 3437 )  100.n
R_D52203LOADxxQSSE13 ( 0 3439 ) COMPLEX( 390., 0.)
R_D52202xxQSSE13 ( 3438 3437 )  100.n
R_D52202LOADxxQSSE13 ( 0 3438 ) COMPLEX( 390., 0.)
R_D52201xxQSSE13 ( 3436 3437 )  100.n
R_D52201LOADxxQSSE13 ( 0 3436 ) COMPLEX( 9.7692,-5.5365)
R_D52103xxQSSE13 ( 3435 3431 )  100.n
R_D52103LOADxxQSSE13 ( 0 3435 ) COMPLEX( 390., 0.)
R_D52102xxQSSE13 ( 3434 3431 )  100.n
R_D52102LOADxxQSSE13 ( 0 3434 ) COMPLEX( 161.6139,-121.2105)
R_D52101xxQSSE13 ( 3433 3431 )  100.n
R_D52101LOADxxQSSE13 ( 0 3433 ) COMPLEX( 390., 0.)
R_D52L1xxQSSE13 ( 0 0 )  1.E+12
R_D52L2xxQSSE13 ( 3429 3437 )  100.n
R_D52307xxQSSE13 ( 3432 3429 )  100.n
R_D52307LOADxxQSSE13 ( 0 3432 ) COMPLEX( 390., 0.)
R_D52104xxQSSE13 ( 3430 3431 )  100.n
R_D52104LOADxxQSSE13 ( 0 3430 ) COMPLEX( 390., 0.)
R_D52308xxQSSE13 ( 3428 3429 )  100.n
R_D52308LOADxxQSSE13 ( 0 3428 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA CCMD3 
R_D52101xxCCMD3 ( 3470 3450 )  100.n
R_D52101LOADxxCCMD3 ( 0 3470 ) COMPLEX( 123.9039,-92.928)
R_D52E1xxCCMD3 ( 479 3450 )  100.n
R_D52209xxCCMD3 ( 3468 3447 )  100.n
R_D52209LOADxxCCMD3 ( 0 3468 ) COMPLEX( 390., 0.)
R_D52E2xxCCMD3 ( 421 3447 )  100.n
R_D52208xxCCMD3 ( 3466 3447 )  100.n
R_D52208LOADxxCCMD3 ( 0 3466 ) COMPLEX( 1.363267K,-1.593835K)
R_D52207xxCCMD3 ( 3465 3447 )  100.n
R_D52207LOADxxCCMD3 ( 0 3465 ) COMPLEX( 235.5726,-188.9955)
R_D52206xxCCMD3 ( 3464 3447 )  100.n
R_D52206LOADxxCCMD3 ( 0 3464 ) COMPLEX( 5.8614,-3.3219)
R_D52205xxCCMD3 ( 3463 3447 )  100.n
R_D52205LOADxxCCMD3 ( 0 3463 ) COMPLEX( 11.6097,-6.8889)
R_D52204xxCCMD3 ( 3462 3447 )  100.n
R_D52204LOADxxCCMD3 ( 0 3462 ) COMPLEX( 390., 0.)
R_D52203xxCCMD3 ( 3461 3447 )  100.n
R_D52203LOADxxCCMD3 ( 0 3461 ) COMPLEX( 1.363267K,-1.593835K)
R_D52202xxCCMD3 ( 3460 3447 )  100.n
R_D52202LOADxxCCMD3 ( 0 3460 ) COMPLEX( 235.5726,-188.9955)
R_D52201xxCCMD3 ( 3459 3447 )  100.n
R_D52201LOADxxCCMD3 ( 0 3459 ) COMPLEX( 123.9039,-92.928)
R_D52110xxCCMD3 ( 3458 3450 )  100.n
R_D52110LOADxxCCMD3 ( 0 3458 ) COMPLEX( 390., 0.)
R_D52109xxCCMD3 ( 3457 3450 )  100.n
R_D52109LOADxxCCMD3 ( 0 3457 ) COMPLEX( 11.6097,-6.8889)
R_D52108xxCCMD3 ( 3456 3450 )  100.n
R_D52108LOADxxCCMD3 ( 0 3456 ) COMPLEX( 11.6097,-6.8889)
R_D52107xxCCMD3 ( 3455 3450 )  100.n
R_D52107LOADxxCCMD3 ( 0 3455 ) COMPLEX( 390., 0.)
R_D52106xxCCMD3 ( 3454 3450 )  100.n
R_D52106LOADxxCCMD3 ( 0 3454 ) COMPLEX( 390., 0.)
R_D52105xxCCMD3 ( 3453 3450 )  100.n
R_D52105LOADxxCCMD3 ( 0 3453 ) COMPLEX( 5.8614,-3.3219)
R_D52104xxCCMD3 ( 3452 3450 )  100.n
R_D52104LOADxxCCMD3 ( 0 3452 ) COMPLEX( 5.8614,-3.3219)
R_D52103xxCCMD3 ( 3451 3450 )  100.n
R_D52103LOADxxCCMD3 ( 0 3451 ) COMPLEX( 390., 0.)
R_D52102xxCCMD3 ( 3449 3450 )  100.n
R_D52102LOADxxCCMD3 ( 0 3449 ) COMPLEX( 1.363267K,-1.593835K)
R_D52LxxCCMD3 ( 0 0 )  1.E+12
R_D52211xxCCMD3 ( 3448 3447 )  100.n
R_D52211LOADxxCCMD3 ( 0 3448 ) COMPLEX( 390., 0.)
R_D52210xxCCMD3 ( 3446 3447 )  100.n
R_D52210LOADxxCCMD3 ( 0 3446 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA CCMD4 
R_D52101xxCCMD4 ( 3495 3475 )  100.n
R_D52101LOADxxCCMD4 ( 0 3495 ) COMPLEX( 123.9039,-92.928)
R_D52E1xxCCMD4 ( 412 3475 )  100.n
R_D52209xxCCMD4 ( 3493 3472 )  100.n
R_D52209LOADxxCCMD4 ( 0 3493 ) COMPLEX( 390., 0.)
R_D52E2xxCCMD4 ( 402 3472 )  100.n
R_D52208xxCCMD4 ( 3491 3472 )  100.n
R_D52208LOADxxCCMD4 ( 0 3491 ) COMPLEX( 1.363267K,-1.593835K)
R_D52207xxCCMD4 ( 3490 3472 )  100.n
R_D52207LOADxxCCMD4 ( 0 3490 ) COMPLEX( 235.5726,-188.9955)
R_D52206xxCCMD4 ( 3489 3472 )  100.n
R_D52206LOADxxCCMD4 ( 0 3489 ) COMPLEX( 5.8614,-3.3219)
R_D52205xxCCMD4 ( 3488 3472 )  100.n
R_D52205LOADxxCCMD4 ( 0 3488 ) COMPLEX( 9.7692,-5.5365)
R_D52204xxCCMD4 ( 3487 3472 )  100.n
R_D52204LOADxxCCMD4 ( 0 3487 ) COMPLEX( 390., 0.)
R_D52203xxCCMD4 ( 3486 3472 )  100.n
R_D52203LOADxxCCMD4 ( 0 3486 ) COMPLEX( 1.363267K,-1.593835K)
R_D52202xxCCMD4 ( 3485 3472 )  100.n
R_D52202LOADxxCCMD4 ( 0 3485 ) COMPLEX( 235.5726,-188.9955)
R_D52201xxCCMD4 ( 3484 3472 )  100.n
R_D52201LOADxxCCMD4 ( 0 3484 ) COMPLEX( 123.9039,-92.928)
R_D52110xxCCMD4 ( 3483 3475 )  100.n
R_D52110LOADxxCCMD4 ( 0 3483 ) COMPLEX( 390., 0.)
R_D52109xxCCMD4 ( 3482 3475 )  100.n
R_D52109LOADxxCCMD4 ( 0 3482 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxCCMD4 ( 3481 3475 )  100.n
R_D52108LOADxxCCMD4 ( 0 3481 ) COMPLEX( 9.7692,-5.5365)
R_D52107xxCCMD4 ( 3480 3475 )  100.n
R_D52107LOADxxCCMD4 ( 0 3480 ) COMPLEX( 390., 0.)
R_D52106xxCCMD4 ( 3479 3475 )  100.n
R_D52106LOADxxCCMD4 ( 0 3479 ) COMPLEX( 390., 0.)
R_D52105xxCCMD4 ( 3478 3475 )  100.n
R_D52105LOADxxCCMD4 ( 0 3478 ) COMPLEX( 5.8614,-3.3219)
R_D52104xxCCMD4 ( 3477 3475 )  100.n
R_D52104LOADxxCCMD4 ( 0 3477 ) COMPLEX( 5.8614,-3.3219)
R_D52103xxCCMD4 ( 3476 3475 )  100.n
R_D52103LOADxxCCMD4 ( 0 3476 ) COMPLEX( 390., 0.)
R_D52102xxCCMD4 ( 3474 3475 )  100.n
R_D52102LOADxxCCMD4 ( 0 3474 ) COMPLEX( 1.363267K,-1.593835K)
R_D52LxxCCMD4 ( 0 0 )  1.E+12
R_D52211xxCCMD4 ( 3473 3472 )  100.n
R_D52211LOADxxCCMD4 ( 0 3473 ) COMPLEX( 390., 0.)
R_D52210xxCCMD4 ( 3471 3472 )  100.n
R_D52210LOADxxCCMD4 ( 0 3471 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA CCME3 
R_D52E1xxCCME3 ( 490 3499 )  100.n
R_D52E2xxCCME3 ( 458 3497 )  100.n
R_D52206xxCCME3 ( 3512 3497 )  100.n
R_D52206LOADxxCCME3 ( 0 3512 ) COMPLEX( 390., 0.)
R_D52205xxCCME3 ( 3511 3497 )  100.n
R_D52205LOADxxCCME3 ( 0 3511 ) COMPLEX( 390., 0.)
R_D52204xxCCME3 ( 3510 3497 )  100.n
R_D52204LOADxxCCME3 ( 0 3510 ) COMPLEX( 26.6742,-17.9253)
R_D52203xxCCME3 ( 3509 3497 )  100.n
R_D52203LOADxxCCME3 ( 0 3509 ) COMPLEX( 390., 0.)
R_D52202xxCCME3 ( 3508 3497 )  100.n
R_D52202LOADxxCCME3 ( 0 3508 ) COMPLEX( 2.8638,-1.6992)
R_D52201xxCCME3 ( 3507 3497 )  100.n
R_D52201LOADxxCCME3 ( 0 3507 ) COMPLEX( 2.8638,-1.6992)
R_D52107xxCCME3 ( 3506 3499 )  100.n
R_D52107LOADxxCCME3 ( 0 3506 ) COMPLEX( 1.363267K,-1.593835K)
R_D52106xxCCME3 ( 3505 3499 )  100.n
R_D52106LOADxxCCME3 ( 0 3505 ) COMPLEX( 390., 0.)
R_D52105xxCCME3 ( 3504 3499 )  100.n
R_D52105LOADxxCCME3 ( 0 3504 ) COMPLEX( 390., 0.)
R_D52104xxCCME3 ( 3503 3499 )  100.n
R_D52104LOADxxCCME3 ( 0 3503 ) COMPLEX( 53.3484,-35.8503)
R_D52103xxCCME3 ( 3502 3499 )  100.n
R_D52103LOADxxCCME3 ( 0 3502 ) COMPLEX( 390., 0.)
R_D52102xxCCME3 ( 3501 3499 )  100.n
R_D52102LOADxxCCME3 ( 0 3501 ) COMPLEX( 2.8638,-1.6992)
R_D52101xxCCME3 ( 3500 3499 )  100.n
R_D52101LOADxxCCME3 ( 0 3500 ) COMPLEX( 2.8638,-1.6992)
R_D52LxxCCME3 ( 0 0 )  1.E+12
R_D52108xxCCME3 ( 3498 3499 )  100.n
R_D52108LOADxxCCME3 ( 0 3498 ) COMPLEX( 390., 0.)
R_D52207xxCCME3 ( 3496 3497 )  100.n
R_D52207LOADxxCCME3 ( 0 3496 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA CCME4 
R_D52E1xxCCME4 ( 407 3516 )  100.n
R_D52E2xxCCME4 ( 400 3514 )  100.n
R_D52206xxCCME4 ( 3529 3514 )  100.n
R_D52206LOADxxCCME4 ( 0 3529 ) COMPLEX( 390., 0.)
R_D52205xxCCME4 ( 3528 3514 )  100.n
R_D52205LOADxxCCME4 ( 0 3528 ) COMPLEX( 390., 0.)
R_D52204xxCCME4 ( 3527 3514 )  100.n
R_D52204LOADxxCCME4 ( 0 3527 ) COMPLEX( 26.6742,-17.9253)
R_D52203xxCCME4 ( 3526 3514 )  100.n
R_D52203LOADxxCCME4 ( 0 3526 ) COMPLEX( 390., 0.)
R_D52202xxCCME4 ( 3525 3514 )  100.n
R_D52202LOADxxCCME4 ( 0 3525 ) COMPLEX( 2.8638,-1.6992)
R_D52201xxCCME4 ( 3524 3514 )  100.n
R_D52201LOADxxCCME4 ( 0 3524 ) COMPLEX( 2.8638,-1.6992)
R_D52107xxCCME4 ( 3523 3516 )  100.n
R_D52107LOADxxCCME4 ( 0 3523 ) COMPLEX( 1.363267K,-1.593835K)
R_D52106xxCCME4 ( 3522 3516 )  100.n
R_D52106LOADxxCCME4 ( 0 3522 ) COMPLEX( 390., 0.)
R_D52105xxCCME4 ( 3521 3516 )  100.n
R_D52105LOADxxCCME4 ( 0 3521 ) COMPLEX( 390., 0.)
R_D52104xxCCME4 ( 3520 3516 )  100.n
R_D52104LOADxxCCME4 ( 0 3520 ) COMPLEX( 53.3484,-35.8503)
R_D52103xxCCME4 ( 3519 3516 )  100.n
R_D52103LOADxxCCME4 ( 0 3519 ) COMPLEX( 390., 0.)
R_D52102xxCCME4 ( 3518 3516 )  100.n
R_D52102LOADxxCCME4 ( 0 3518 ) COMPLEX( 2.8638,-1.6992)
R_D52101xxCCME4 ( 3517 3516 )  100.n
R_D52101LOADxxCCME4 ( 0 3517 ) COMPLEX( 2.8638,-1.6992)
R_D52LxxCCME4 ( 0 0 )  1.E+12
R_D52108xxCCME4 ( 3515 3516 )  100.n
R_D52108LOADxxCCME4 ( 0 3515 ) COMPLEX( 390., 0.)
R_D52207xxCCME4 ( 3513 3514 )  100.n
R_D52207LOADxxCCME4 ( 0 3513 ) COMPLEX( 390., 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSAM3 
R_D52101xxQSAM3 ( 3531 3561 )  100.n
R_D52101LOADxxQSAM3 ( 0 3561 ) COMPLEX( 21.6276,-14.5338)
R_D52102xxQSAM3 ( 3560 3531 )  100.n
R_D52102LOADxxQSAM3 ( 0 3560 ) COMPLEX( 390., 0.)
R_D52103xxQSAM3 ( 3559 3531 )  100.n
R_D52103LOADxxQSAM3 ( 0 3559 ) COMPLEX( 86.7843,-60.576)
R_D52104xxQSAM3 ( 3558 3531 )  100.n
R_D52104LOADxxQSAM3 ( 0 3558 ) COMPLEX( 168.96,-126.72)
R_D52105xxQSAM3 ( 3557 3531 )  100.n
R_D52105LOADxxQSAM3 ( 0 3557 ) COMPLEX( 390., 0.)
R_D52106xxQSAM3 ( 3556 3531 )  100.n
R_D52106LOADxxQSAM3 ( 0 3556 ) COMPLEX( 21.6276,-14.5338)
R_D52107LOADxxQSAM3 ( 0 3555 ) COMPLEX( 21.6276,-14.5338)
R_D52107xxQSAM3 ( 3555 3531 )  100.n
R_D52109xxQSAM3 ( 3554 3531 )  100.n
R_D52109LOADxxQSAM3 ( 3554 0 ) COMPLEX( 390., 0.)
R_D52110xxQSAM3 ( 3553 3531 )  100.n
R_D52110LOADxxQSAM3 ( 3553 0 ) COMPLEX( 71.0055,-49.5621)
R_D52111xxQSAM3 ( 3552 3531 )  100.n
R_D52111LOADxxQSAM3 ( 3552 0 ) COMPLEX( 390., 0.)
R_D52112xxQSAM3 ( 3551 3531 )  100.n
R_D52112LOADxxQSAM3 ( 3551 0 ) COMPLEX( 5.8614,-3.3219)
R_D52113xxQSAM3 ( 3550 3531 )  100.n
R_D52113LOADxxQSAM3 ( 3550 0 ) COMPLEX( 21.6276,-14.5338)
R_D52114xxQSAM3 ( 3549 3531 )  100.n
R_D52114LOADxxQSAM3 ( 3549 0 ) COMPLEX( 53.3484,-35.8503)
R_D52ExxQSAM3 ( 602 3531 )  100.n
R_D52115xxQSAM3 ( 3547 3531 )  100.n
R_D52115LOADxxQSAM3 ( 3547 0 ) COMPLEX( 390., 0.)
R_D52117xxQSAM3 ( 3531 3546 )  100.n
R_D52117LOADxxQSAM3 ( 0 3546 ) COMPLEX( 39.204,-18.9873)
R_D52118xxQSAM3 ( 3545 3531 )  100.n
R_D52118LOADxxQSAM3 ( 0 3545 ) COMPLEX( 25.998,-11.8449)
R_D52119xxQSAM3 ( 3544 3531 )  100.n
R_D52119LOADxxQSAM3 ( 0 3544 ) COMPLEX( 390., 0.)
R_D52120xxQSAM3 ( 3543 3531 )  100.n
R_D52120LOADxxQSAM3 ( 0 3543 ) COMPLEX( 7.7439, 0.)
R_D52121xxQSAM3 ( 3542 3531 )  100.n
R_D52121LOADxxQSAM3 ( 0 3542 ) COMPLEX( 355.0272,-247.8105)
R_D52122xxQSAM3 ( 3541 3531 )  100.n
R_D52122LOADxxQSAM3 ( 0 3541 ) COMPLEX( 390., 0.)
R_D52116LOADxxQSAM3 ( 0 3540 ) COMPLEX( 39.204,-18.9873)
R_D52116xxQSAM3 ( 3540 3531 )  100.n
R_D52123xxQSAM3 ( 3539 3531 )  100.n
R_D52123LOADxxQSAM3 ( 3539 0 ) COMPLEX( 4.6578,-2.256)
R_D52124xxQSAM3 ( 3538 3531 )  100.n
R_D52124LOADxxQSAM3 ( 3538 0 ) COMPLEX( 390., 0.)
R_D52125xxQSAM3 ( 3537 3531 )  100.n
R_D52125LOADxxQSAM3 ( 3537 0 ) COMPLEX( 2.4516,-0.8058)
R_D52126xxQSAM3 ( 3536 3531 )  100.n
R_D52126LOADxxQSAM3 ( 3536 0 ) COMPLEX( 390., 0.)
R_D52127xxQSAM3 ( 3535 3531 )  100.n
R_D52127LOADxxQSAM3 ( 3535 0 ) COMPLEX( 2.6571,-1.1319)
R_D52128xxQSAM3 ( 3534 3531 )  100.n
R_D52128LOADxxQSAM3 ( 3534 0 ) COMPLEX( 1.3287,-0.5661)
R_D52129xxQSAM3 ( 3533 3531 )  100.n
R_D52129LOADxxQSAM3 ( 3533 0 ) COMPLEX( 1.8498,-0.8427)
R_D52130xxQSAM3 ( 3532 3531 )  100.n
R_D52130LOADxxQSAM3 ( 3532 0 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSAM3 ( 0 3530 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxQSAM3 ( 3530 3531 )  100.n
*----------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Aux CA QSAM4 
R_D52101xxQSAM4 ( 3563 3593 )  100.n
R_D52101LOADxxQSAM4 ( 0 3593 ) COMPLEX( 21.6276,-14.5338)
R_D52102xxQSAM4 ( 3592 3563 )  100.n
R_D52102LOADxxQSAM4 ( 0 3592 ) COMPLEX( 390., 0.)
R_D52103xxQSAM4 ( 3591 3563 )  100.n
R_D52103LOADxxQSAM4 ( 0 3591 ) COMPLEX( 86.7843,-60.576)
R_D52104xxQSAM4 ( 3590 3563 )  100.n
R_D52104LOADxxQSAM4 ( 0 3590 ) COMPLEX( 168.96,-126.72)
R_D52105xxQSAM4 ( 3589 3563 )  100.n
R_D52105LOADxxQSAM4 ( 0 3589 ) COMPLEX( 390., 0.)
R_D52106xxQSAM4 ( 3588 3563 )  100.n
R_D52106LOADxxQSAM4 ( 0 3588 ) COMPLEX( 21.6276,-14.5338)
R_D52107LOADxxQSAM4 ( 0 3587 ) COMPLEX( 21.6276,-14.5338)
R_D52107xxQSAM4 ( 3587 3563 )  100.n
R_D52109xxQSAM4 ( 3586 3563 )  100.n
R_D52109LOADxxQSAM4 ( 3586 0 ) COMPLEX( 390., 0.)
R_D52110xxQSAM4 ( 3585 3563 )  100.n
R_D52110LOADxxQSAM4 ( 3585 0 ) COMPLEX( 71.0055,-49.5621)
R_D52111xxQSAM4 ( 3584 3563 )  100.n
R_D52111LOADxxQSAM4 ( 3584 0 ) COMPLEX( 390., 0.)
R_D52112xxQSAM4 ( 3583 3563 )  100.n
R_D52112LOADxxQSAM4 ( 3583 0 ) COMPLEX( 5.8614,-3.3219)
R_D52113xxQSAM4 ( 3582 3563 )  100.n
R_D52113LOADxxQSAM4 ( 3582 0 ) COMPLEX( 21.6276,-14.5338)
R_D52114xxQSAM4 ( 3581 3563 )  100.n
R_D52114LOADxxQSAM4 ( 3581 0 ) COMPLEX( 53.3484,-35.8503)
R_D52ExxQSAM4 ( 533 3563 )  100.n
R_D52115xxQSAM4 ( 3579 3563 )  100.n
R_D52115LOADxxQSAM4 ( 3579 0 ) COMPLEX( 390., 0.)
R_D52117xxQSAM4 ( 3563 3578 )  100.n
R_D52117LOADxxQSAM4 ( 0 3578 ) COMPLEX( 39.204,-18.9873)
R_D52118xxQSAM4 ( 3577 3563 )  100.n
R_D52118LOADxxQSAM4 ( 0 3577 ) COMPLEX( 25.998,-11.8449)
R_D52119xxQSAM4 ( 3576 3563 )  100.n
R_D52119LOADxxQSAM4 ( 0 3576 ) COMPLEX( 390., 0.)
R_D52120xxQSAM4 ( 3575 3563 )  100.n
R_D52120LOADxxQSAM4 ( 0 3575 ) COMPLEX( 7.7439, 0.)
R_D52121xxQSAM4 ( 3574 3563 )  100.n
R_D52121LOADxxQSAM4 ( 0 3574 ) COMPLEX( 355.0272,-247.8105)
R_D52122xxQSAM4 ( 3573 3563 )  100.n
R_D52122LOADxxQSAM4 ( 0 3573 ) COMPLEX( 390., 0.)
R_D52116LOADxxQSAM4 ( 0 3572 ) COMPLEX( 39.204,-18.9873)
R_D52116xxQSAM4 ( 3572 3563 )  100.n
R_D52123xxQSAM4 ( 3571 3563 )  100.n
R_D52123LOADxxQSAM4 ( 3571 0 ) COMPLEX( 4.6578,-2.256)
R_D52124xxQSAM4 ( 3570 3563 )  100.n
R_D52124LOADxxQSAM4 ( 3570 0 ) COMPLEX( 390., 0.)
R_D52125xxQSAM4 ( 3569 3563 )  100.n
R_D52125LOADxxQSAM4 ( 3569 0 ) COMPLEX( 2.4516,-0.8058)
R_D52126xxQSAM4 ( 3568 3563 )  100.n
R_D52126LOADxxQSAM4 ( 3568 0 ) COMPLEX( 390., 0.)
R_D52127xxQSAM4 ( 3567 3563 )  100.n
R_D52127LOADxxQSAM4 ( 3567 0 ) COMPLEX( 2.6571,-1.1319)
R_D52128xxQSAM4 ( 3566 3563 )  100.n
R_D52128LOADxxQSAM4 ( 3566 0 ) COMPLEX( 1.3287,-0.5661)
R_D52129xxQSAM4 ( 3565 3563 )  100.n
R_D52129LOADxxQSAM4 ( 3565 0 ) COMPLEX( 1.8498,-0.8427)
R_D52130xxQSAM4 ( 3564 3563 )  100.n
R_D52130LOADxxQSAM4 ( 3564 0 ) COMPLEX( 390., 0.)
R_D52108LOADxxQSAM4 ( 0 3562 ) COMPLEX( 9.7692,-5.5365)
R_D52108xxQSAM4 ( 3562 3563 )  100.n
