TITLE UH JIRAU POWER FLOW (March/2018) 
* -------------------------------------------------------------------------------- 
* Notes: 
* TO-DO1: capacitors in shunt mode to the circuit breaker. 
* TO-DO2: ... 
* TO-DO3: ... 
* -------------------------------------------------------------------------------- 
* Models 
* A magnetic coupling 13.8kV to 525kV: 
.subckt COUPLING_525K  ( 1 3 )
*1,2: primary nodes 
*2,3: secondary nodes 
*13.8kV to 525kV 
Lsecondary ( 0 3 )  2.894612K
Lprimary ( 0 1 )  2.
K  Lsecondary  Lprimary  0.9999999
.ends COUPLING_525K
* 
*Version 3: 2 independent monophasic transformers in parallel. 
.subckt MONOPHASIC_TRANSFORMER_525K  ( 1 2 3 )
*1,0: primary A 
*2,0: primary B 
*3,0: secondary 
XTEa ( 1 3 )  COUPLING_525K
XTEb ( 2 3 )  COUPLING_525K
.ends MONOPHASIC_TRANSFORMER_525K
* 
* A magnetic coupling 13.8kV to 440V: 
.subckt MONOPHASIC_TRANSFORMER_440  ( 1 2 )
*1,0: primary nodes 
*2,0: secondary nodes 
*13.8kV to 440V 
Lsecondary ( 0 2 )  2.033186
Lprimary ( 0 1 )  2.K
K  Lsecondary  Lprimary  0.9999999
.ends MONOPHASIC_TRANSFORMER_440
* 
* A magnetic coupling where a=1: 
.subckt MONOPHASIC_REGULATOR  ( 1 2 )
*1,0: primary nodes 
*2,0: secondary nodes 
*a=1 
Lsecondary ( 0 2 )  2.K
Lprimary ( 0 1 )  2.K
K  Lsecondary  Lprimary  0.9999999
.ends MONOPHASIC_REGULATOR
* 
* LT1 and LT2: 
.subckt LT_LT1_LT2  ( 1 2 )
***R_LT1_PI ( 1 2 ) COMPLEX( 1.624, 28.765) 
R_LT1_PI ( 1 2 ) COMPLEX( 1.624, 0.)
***R_LT1_PI1 ( 1 0 ) COMPLEX( 0.,-4.05351K) 
***R_LT1_PI2 ( 2 0 ) COMPLEX( 0.,-4.05351K) 
.ends LT_LT1_LT2
* LT3: 
.subckt LT_LT3  ( 1 2 )
***R_LT3_PI ( 1 2 ) COMPLEX( 32.344, 122.882) 
R_LT3_PI ( 1 2 ) COMPLEX( 1.624, 0.)
.ends LT_LT3
* LT4 and LT5: 
.subckt LT_LT45  ( 1 2 )
***R_LT45_PI ( 1 2 ) COMPLEX( 1.624, 0.) 
R_LT45_PI ( 1 2 ) COMPLEX( 100.n, 0.)
.ends LT_LT45
* 
* 
* -------------------------------------------------------------------------------- 
* Netlist: SE MD, SE ME and SE Coletora 

R_D52A1_5 ( 175 176 ) COMPLEX( 100.n, 0.)
R_D52A1_6 ( 166 167 ) COMPLEX( 100.n, 0.)
R_D52BT_1 ( 65 179 ) COMPLEX( 100.n, 0.)
R_D52BT_2 ( 59 181 ) COMPLEX( 100.n, 0.)
R_D52C1_4 ( 168 163 ) COMPLEX( 100.n, 0.)
R_D52C1_5 ( 173 172 ) COMPLEX( 100.n, 0.)
R_D52C1_6 ( 164 162 ) COMPLEX( 100.n, 0.)
R_D52G_1 ( 110 229 ) COMPLEX( 100.n, 0.)
R_D52G_10 ( 115 235 ) COMPLEX( 100.n, 0.)
R_D52G_11 ( 113 236 ) COMPLEX( 100.n, 0.)
R_D52G_12 ( 112 237 ) COMPLEX( 100.n, 0.)
R_D52G_13 ( 122 238 ) COMPLEX( 100.n, 0.)
R_D52G_14 ( 121 239 ) COMPLEX( 100.n, 0.)
R_D52G_15 ( 119 240 ) COMPLEX( 100.n, 0.)
R_D52G_16 ( 118 241 ) COMPLEX( 100.n, 0.)
R_D52G_17 ( 128 223 ) COMPLEX( 100.n, 0.)
R_D52G_18 ( 127 224 ) COMPLEX( 100.n, 0.)
R_D52G_19 ( 125 225 ) COMPLEX( 100.n, 0.)
R_D52G_2 ( 109 228 ) COMPLEX( 100.n, 0.)
R_D52G_20 ( 124 222 ) COMPLEX( 100.n, 0.)
R_D52G_21 ( 200 134 ) COMPLEX( 100.n, 0.)
R_D52G_22 ( 133 201 ) COMPLEX( 100.n, 0.)
R_D52G_23 ( 202 131 ) COMPLEX( 100.n, 0.)
R_D52G_24 ( 130 203 ) COMPLEX( 100.n, 0.)
R_D52G_25 ( 140 196 ) COMPLEX( 100.n, 0.)
R_D52G_26 ( 139 197 ) COMPLEX( 100.n, 0.)
R_D52G_27 ( 137 198 ) COMPLEX( 100.n, 0.)
R_D52G_28 ( 136 199 ) COMPLEX( 100.n, 0.)
R_D52G_29 ( 221 158 ) COMPLEX( 100.n, 0.)
R_D52G_3 ( 107 227 ) COMPLEX( 100.n, 0.)
R_D52G_30 ( 220 157 ) COMPLEX( 100.n, 0.)
R_D52G_31 ( 155 219 ) COMPLEX( 100.n, 0.)
R_D52G_32 ( 218 154 ) COMPLEX( 100.n, 0.)
R_D52G_33 ( 217 152 ) COMPLEX( 100.n, 0.)
R_D52G_34 ( 216 151 ) COMPLEX( 100.n, 0.)
R_D52G_35 ( 215 149 ) COMPLEX( 100.n, 0.)
R_D52G_36 ( 214 148 ) COMPLEX( 100.n, 0.)
R_D52G_37 ( 146 213 ) COMPLEX( 100.n, 0.)
R_D52G_38 ( 212 145 ) COMPLEX( 100.n, 0.)
R_D52G_39 ( 143 211 ) COMPLEX( 100.n, 0.)
R_D52G_4 ( 106 226 ) COMPLEX( 100.n, 0.)
R_D52G_40 ( 210 142 ) COMPLEX( 100.n, 0.)
R_D52G_41 ( 192 98 ) COMPLEX( 100.n, 0.)
R_D52G_42 ( 97 193 ) COMPLEX( 100.n, 0.)
R_D52G_43 ( 194 95 ) COMPLEX( 100.n, 0.)
R_D52G_44 ( 94 195 ) COMPLEX( 100.n, 0.)
R_D52G_45 ( 92 209 ) COMPLEX( 100.n, 0.)
R_D52G_46 ( 208 91 ) COMPLEX( 100.n, 0.)
R_D52G_47 ( 89 207 ) COMPLEX( 100.n, 0.)
R_D52G_48 ( 206 88 ) COMPLEX( 100.n, 0.)
R_D52G_49 ( 86 205 ) COMPLEX( 100.n, 0.)
R_D52G_5 ( 104 233 ) COMPLEX( 100.n, 0.)
R_D52G_50 ( 84 204 ) COMPLEX( 100.n, 0.)
R_D52G_6 ( 103 232 ) COMPLEX( 100.n, 0.)
R_D52G_7 ( 101 231 ) COMPLEX( 100.n, 0.)
R_D52G_8 ( 100 230 ) COMPLEX( 100.n, 0.)
R_D52G_9 ( 116 234 ) COMPLEX( 100.n, 0.)
R_D52L_1 ( 72 186 ) COMPLEX( 100.n, 0.)
R_D52L_2 ( 64 185 ) COMPLEX( 100.n, 0.)
R_D52L_3 ( 57 184 ) COMPLEX( 100.n, 0.)
R_D52L_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L_5 ( 60 188 ) COMPLEX( 100.n, 0.)
R_D52RE0_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52T_1 ( 243 70 ) COMPLEX( 100.n, 0.)
R_D52T_10 ( 78 252 ) COMPLEX( 100.n, 0.)
R_D52T_11 ( 251 82 ) COMPLEX( 100.n, 0.)
R_D52T_12 ( 248 159 ) COMPLEX( 100.n, 0.)
R_D52T_13 ( 160 246 ) COMPLEX( 100.n, 0.)
R_D52T_2 ( 245 71 ) COMPLEX( 100.n, 0.)
R_D52T_3 ( 267 68 ) COMPLEX( 100.n, 0.)
R_D52T_4 ( 264 67 ) COMPLEX( 100.n, 0.)
R_D52T_5 ( 262 74 ) COMPLEX( 100.n, 0.)
R_D52T_6 ( 75 261 ) COMPLEX( 100.n, 0.)
R_D52T_7 ( 258 76 ) COMPLEX( 100.n, 0.)
R_D52T_8 ( 256 80 ) COMPLEX( 100.n, 0.)
R_D52T_9 ( 79 254 ) COMPLEX( 100.n, 0.)
R_S57B1_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B1_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B2_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B2_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B3_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B3_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B4_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57B4_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57BT1_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57BT1_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57BT2_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57BT2_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L1_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L1_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L1_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L1_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L1_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L2_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L2_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L2_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L2_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L2_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L3_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L3_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L3_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L3_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57L3_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57LA1_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57LA1_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57LA1_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T1_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T2_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57T3_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_14 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_15 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_16 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_17 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_18 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_19 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_20 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_21 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_22 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_23 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_24 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_25 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_26 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_27 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_28 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_29 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_30 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_31 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_32 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_33 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_34 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_35 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_36 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_37 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_38 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_39 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_40 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_41 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_42 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_43 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_44 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_45 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_46 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_47 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_48 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_49 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_50 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TA_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_14 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_15 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_16 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_17 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_18 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_19 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_20 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_21 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_22 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_23 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_24 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_25 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_26 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_27 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_28 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_29 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_30 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_31 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_32 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_33 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_34 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_35 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_36 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_37 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_38 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_39 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_40 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_41 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_42 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_43 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_44 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_45 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_46 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_47 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_48 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_49 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_50 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S57TB_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89A1_4 ( 171 51 ) COMPLEX( 100.n, 0.)
R_S89A1_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89A1_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89AC1_4 ( 169 170 ) COMPLEX( 100.n, 0.)
R_S89AC1_5 ( 174 175 ) COMPLEX( 100.n, 0.)
R_S89AC1_6 ( 165 166 ) COMPLEX( 100.n, 0.)
R_S89B1_1 ( 63 180 ) COMPLEX( 100.n, 0.)
R_S89B1_2 ( 190 69 ) COMPLEX( 100.n, 0.)
R_S89B2_1 ( 180 191 ) COMPLEX( 100.n, 0.)
R_S89B2_2 ( 66 190 ) COMPLEX( 100.n, 0.)
R_S89B3_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89B3_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89B4_1 ( 56 182 ) COMPLEX( 100.n, 0.)
R_S89B4_2 ( 178 183 ) COMPLEX( 100.n, 0.)
R_S89B5_1 ( 56 177 ) COMPLEX( 100.n, 0.)
R_S89B5_2 ( 81 178 ) COMPLEX( 100.n, 0.)
R_S89B6_1 ( 61 191 ) COMPLEX( 100.n, 0.)
R_S89B6_2 ( 73 66 ) COMPLEX( 100.n, 0.)
R_S89BTA_1 ( 179 180 ) COMPLEX( 100.n, 0.)
R_S89BTA_2 ( 181 182 ) COMPLEX( 100.n, 0.)
R_S89BTB_1 ( 65 190 ) COMPLEX( 100.n, 0.)
R_S89BTB_2 ( 59 183 ) COMPLEX( 100.n, 0.)
R_S89CA1_4 ( 168 169 ) COMPLEX( 100.n, 0.)
R_S89CA1_5 ( 173 174 ) COMPLEX( 100.n, 0.)
R_S89CA1_6 ( 164 165 ) COMPLEX( 100.n, 0.)
R_S89CB1_4 ( 163 50 ) COMPLEX( 100.n, 0.)
R_S89CB1_5 ( 50 172 ) COMPLEX( 100.n, 0.)
R_S89CB1_6 ( 162 50 ) COMPLEX( 100.n, 0.)
R_S89G_1 ( 229 108 ) COMPLEX( 100.n, 0.)
R_S89G_10 ( 235 114 ) COMPLEX( 100.n, 0.)
R_S89G_11 ( 236 111 ) COMPLEX( 100.n, 0.)
R_S89G_12 ( 237 111 ) COMPLEX( 100.n, 0.)
R_S89G_13 ( 238 120 ) COMPLEX( 100.n, 0.)
R_S89G_14 ( 239 120 ) COMPLEX( 100.n, 0.)
R_S89G_15 ( 240 117 ) COMPLEX( 100.n, 0.)
R_S89G_16 ( 241 117 ) COMPLEX( 100.n, 0.)
R_S89G_17 ( 223 126 ) COMPLEX( 100.n, 0.)
R_S89G_18 ( 224 126 ) COMPLEX( 100.n, 0.)
R_S89G_19 ( 225 123 ) COMPLEX( 100.n, 0.)
R_S89G_2 ( 228 108 ) COMPLEX( 100.n, 0.)
R_S89G_20 ( 222 123 ) COMPLEX( 100.n, 0.)
R_S89G_21 ( 132 200 ) COMPLEX( 100.n, 0.)
R_S89G_22 ( 201 132 ) COMPLEX( 100.n, 0.)
R_S89G_23 ( 129 202 ) COMPLEX( 100.n, 0.)
R_S89G_24 ( 129 203 ) COMPLEX( 100.n, 0.)
R_S89G_25 ( 196 138 ) COMPLEX( 100.n, 0.)
R_S89G_26 ( 197 138 ) COMPLEX( 100.n, 0.)
R_S89G_27 ( 198 135 ) COMPLEX( 100.n, 0.)
R_S89G_28 ( 199 135 ) COMPLEX( 100.n, 0.)
R_S89G_29 ( 156 221 ) COMPLEX( 100.n, 0.)
R_S89G_3 ( 227 105 ) COMPLEX( 100.n, 0.)
R_S89G_30 ( 156 220 ) COMPLEX( 100.n, 0.)
R_S89G_31 ( 219 153 ) COMPLEX( 100.n, 0.)
R_S89G_32 ( 153 218 ) COMPLEX( 100.n, 0.)
R_S89G_33 ( 150 217 ) COMPLEX( 100.n, 0.)
R_S89G_34 ( 150 216 ) COMPLEX( 100.n, 0.)
R_S89G_35 ( 147 215 ) COMPLEX( 100.n, 0.)
R_S89G_36 ( 147 214 ) COMPLEX( 100.n, 0.)
R_S89G_37 ( 213 144 ) COMPLEX( 100.n, 0.)
R_S89G_38 ( 144 212 ) COMPLEX( 100.n, 0.)
R_S89G_39 ( 211 141 ) COMPLEX( 100.n, 0.)
R_S89G_4 ( 226 105 ) COMPLEX( 100.n, 0.)
R_S89G_40 ( 141 210 ) COMPLEX( 100.n, 0.)
R_S89G_41 ( 96 192 ) COMPLEX( 100.n, 0.)
R_S89G_42 ( 193 96 ) COMPLEX( 100.n, 0.)
R_S89G_43 ( 93 194 ) COMPLEX( 100.n, 0.)
R_S89G_44 ( 93 195 ) COMPLEX( 100.n, 0.)
R_S89G_45 ( 209 90 ) COMPLEX( 100.n, 0.)
R_S89G_46 ( 90 208 ) COMPLEX( 100.n, 0.)
R_S89G_47 ( 207 87 ) COMPLEX( 100.n, 0.)
R_S89G_48 ( 87 206 ) COMPLEX( 100.n, 0.)
R_S89G_49 ( 205 85 ) COMPLEX( 100.n, 0.)
R_S89G_5 ( 233 102 ) COMPLEX( 100.n, 0.)
R_S89G_50 ( 83 204 ) COMPLEX( 100.n, 0.)
R_S89G_6 ( 232 102 ) COMPLEX( 100.n, 0.)
R_S89G_7 ( 231 99 ) COMPLEX( 100.n, 0.)
R_S89G_8 ( 230 99 ) COMPLEX( 100.n, 0.)
R_S89G_9 ( 234 114 ) COMPLEX( 100.n, 0.)
R_S89LA_1 ( 72 63 ) COMPLEX( 100.n, 0.)
R_S89LA_2 ( 64 63 ) COMPLEX( 100.n, 0.)
R_S89LA_3 ( 56 57 ) COMPLEX( 100.n, 0.)
R_S89LA_4 ( 62 61 ) COMPLEX( 100.n, 0.)
R_S89LA_5 ( 60 58 ) COMPLEX( 100.n, 0.)
R_S89LA1_4 ( 269 169 ) COMPLEX( 100.n, 0.)
R_S89LA1_5 ( 270 174 ) COMPLEX( 100.n, 0.)
R_S89LA1_6 ( 268 165 ) COMPLEX( 100.n, 0.)
R_S89LB_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89LB_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89LB_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89LB_4 ( 62 73 ) COMPLEX( 100.n, 0.)
R_S89LB_5 ( 60 77 ) COMPLEX( 100.n, 0.)
R_S89LC_1 ( 53 186 ) COMPLEX( 100.n, 0.)
R_S89LC_2 ( 54 185 ) COMPLEX( 100.n, 0.)
R_S89LC_3 ( 52 184 ) COMPLEX( 100.n, 0.)
R_S89LC_4 ( 187 189 ) COMPLEX( 100.n, 0.)
R_S89LC_5 ( 3594 188 ) COMPLEX( 100.n, 0.)
R_S89LE_1 ( 53 63 ) COMPLEX( 100.n, 0.)
R_S89LE_2 ( 54 63 ) COMPLEX( 100.n, 0.)
R_S89LE_3 ( 56 52 ) COMPLEX( 100.n, 0.)
R_S89LE_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89LE_5 ( 3594 58 ) COMPLEX( 100.n, 0.)
R_S89RE1_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89RE1_5 ( 270 55 ) COMPLEX( 100.n, 0.)
R_S89RE1_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TA_9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S89TB_1 ( 70 69 ) COMPLEX( 100.n, 0.)
R_S89TB_10 ( 77 78 ) COMPLEX( 100.n, 0.)
R_S89TB_11 ( 81 82 ) COMPLEX( 100.n, 0.)
R_S89TB_12 ( 81 159 ) COMPLEX( 100.n, 0.)
R_S89TB_13 ( 81 160 ) COMPLEX( 100.n, 0.)
R_S89TB_2 ( 71 69 ) COMPLEX( 100.n, 0.)
R_S89TB_3 ( 68 66 ) COMPLEX( 100.n, 0.)
R_S89TB_4 ( 67 66 ) COMPLEX( 100.n, 0.)
R_S89TB_5 ( 74 73 ) COMPLEX( 100.n, 0.)
R_S89TB_6 ( 75 73 ) COMPLEX( 100.n, 0.)
R_S89TB_7 ( 76 73 ) COMPLEX( 100.n, 0.)
R_S89TB_8 ( 77 80 ) COMPLEX( 100.n, 0.)
R_S89TB_9 ( 77 79 ) COMPLEX( 100.n, 0.)
R_S89TC_1 ( 243 242 ) COMPLEX( 100.n, 0.)
R_S89TC_10 ( 252 253 ) COMPLEX( 100.n, 0.)
R_S89TC_11 ( 251 250 ) COMPLEX( 100.n, 0.)
R_S89TC_12 ( 248 249 ) COMPLEX( 100.n, 0.)
R_S89TC_13 ( 246 247 ) COMPLEX( 100.n, 0.)
R_S89TC_2 ( 245 244 ) COMPLEX( 100.n, 0.)
R_S89TC_3 ( 267 266 ) COMPLEX( 100.n, 0.)
R_S89TC_4 ( 264 265 ) COMPLEX( 100.n, 0.)
R_S89TC_5 ( 262 263 ) COMPLEX( 100.n, 0.)
R_S89TC_6 ( 261 260 ) COMPLEX( 100.n, 0.)
R_S89TC_7 ( 258 259 ) COMPLEX( 100.n, 0.)
R_S89TC_8 ( 256 257 ) COMPLEX( 100.n, 0.)
R_S89TC_9 ( 254 255 ) COMPLEX( 100.n, 0.)
***R_LT45_METER ( 3594 187 ) COMPLEX( 100.n , 0.) 
X_LT45 ( 3602 3601 )  LT_LT45
R_LT45_METER ( 187 3601 ) COMPLEX( 100.n, 0.)
R_LT45_METER1 ( 3594 3602 ) COMPLEX( 100.n, 0.)
****** 
* Internal current source resistance: 
R_UG01 ( 0 8 ) COMPLEX( 100.n, 0.)
R_UG02 ( 0 7 ) COMPLEX( 100.n, 0.)
R_UG03 ( 0 9 ) COMPLEX( 100.n, 0.)
R_UG04 ( 0 6 ) COMPLEX( 100.n, 0.)
****** 
* Internal voltage source resistance: 
R_UG05 ( 0 4 ) COMPLEX( 100.n, 0.)
R_UG06 ( 0 3 ) COMPLEX( 100.n, 0.)
R_UG07 ( 0 5 ) COMPLEX( 100.n, 0.)
R_UG08 ( 0 2 ) COMPLEX( 100.n, 0.)
R_UG09 ( 0 12 ) COMPLEX( 100.n, 0.)
R_UG10 ( 0 11 ) COMPLEX( 100.n, 0.)
R_UG11 ( 0 13 ) COMPLEX( 100.n, 0.)
R_UG12 ( 0 10 ) COMPLEX( 100.n, 0.)
R_UG13 ( 0 16 ) COMPLEX( 100.n, 0.)
R_UG14 ( 0 15 ) COMPLEX( 100.n, 0.)
R_UG15 ( 0 17 ) COMPLEX( 100.n, 0.)
R_UG16 ( 0 14 ) COMPLEX( 100.n, 0.)
R_UG17 ( 0 20 ) COMPLEX( 100.n, 0.)
R_UG18 ( 0 19 ) COMPLEX( 100.n, 0.)
R_UG19 ( 0 21 ) COMPLEX( 100.n, 0.)
R_UG20 ( 0 18 ) COMPLEX( 100.n, 0.)
R_UG21 ( 0 24 ) COMPLEX( 100.n, 0.)
R_UG22 ( 0 23 ) COMPLEX( 100.n, 0.)
R_UG23 ( 0 25 ) COMPLEX( 100.n, 0.)
R_UG24 ( 0 22 ) COMPLEX( 100.n, 0.)
R_UG25 ( 0 28 ) COMPLEX( 100.n, 0.)
R_UG26 ( 0 27 ) COMPLEX( 100.n, 0.)
R_UG27 ( 0 29 ) COMPLEX( 100.n, 0.)
R_UG28 ( 0 26 ) COMPLEX( 100.n, 0.)
R_UG29 ( 0 32 ) COMPLEX( 100.n, 0.)
R_UG30 ( 0 31 ) COMPLEX( 100.n, 0.)
R_UG31 ( 0 33 ) COMPLEX( 100.n, 0.)
R_UG32 ( 0 30 ) COMPLEX( 100.n, 0.)
R_UG33 ( 0 36 ) COMPLEX( 100.n, 0.)
R_UG34 ( 0 35 ) COMPLEX( 100.n, 0.)
R_UG35 ( 0 37 ) COMPLEX( 100.n, 0.)
R_UG36 ( 0 34 ) COMPLEX( 100.n, 0.)
R_UG37 ( 0 40 ) COMPLEX( 100.n, 0.)
R_UG38 ( 0 39 ) COMPLEX( 100.n, 0.)
R_UG39 ( 0 41 ) COMPLEX( 100.n, 0.)
R_UG40 ( 0 38 ) COMPLEX( 100.n, 0.)
R_UG41 ( 0 44 ) COMPLEX( 100.n, 0.)
R_UG42 ( 0 43 ) COMPLEX( 100.n, 0.)
R_UG43 ( 0 45 ) COMPLEX( 100.n, 0.)
R_UG44 ( 0 42 ) COMPLEX( 100.n, 0.)
R_UG45 ( 0 48 ) COMPLEX( 100.n, 0.)
R_UG46 ( 0 47 ) COMPLEX( 100.n, 0.)
R_UG47 ( 0 49 ) COMPLEX( 100.n, 0.)
R_UG48 ( 0 46 ) COMPLEX( 100.n, 0.)
R_UG49 ( 0 161 ) COMPLEX( 100.n, 0.)
R_UG50 ( 0 1 ) COMPLEX( 100.n, 0.)
**** Valor da resistência no modo fonte de tensão 0.214245 
* For infinite bar load: 
****I_UG01 ( 110 8 ) COMPLEX( 1.0K, 0.) 
****I_UG02 ( 109 7 ) COMPLEX( 1.0K, 0.) 
I_UG01 ( 8 110 ) COMPLEX( 10.0409K, 0.)
I_UG02 ( 7 109 ) COMPLEX( 10.0409K, 7.53066K)
I_UG03 ( 9 107 ) COMPLEX( 10.0409K, 7.53066K)
I_UG04 ( 6 106 ) COMPLEX( 10.0409K, 7.53066K)
I_UG05 ( 4 104 ) COMPLEX( 7.53066K, 0.)
I_UG06 ( 3 103 ) COMPLEX( 7.53066K, 0.)
I_UG07 ( 5 101 ) COMPLEX( 7.53066K, 0.)
I_UG08 ( 2 100 ) COMPLEX( 7.53066K, 0.)
I_UG09 ( 12 116 ) COMPLEX( 7.53066K, 0.)
I_UG10 ( 11 115 ) COMPLEX( 7.53066K, 0.)
I_UG11 ( 13 113 ) COMPLEX( 7.53066K, 0.)
I_UG12 ( 10 112 ) COMPLEX( 7.53066K, 0.)
I_UG13 ( 16 122 ) COMPLEX( 7.53066K, 0.)
I_UG14 ( 15 121 ) COMPLEX( 7.53066K, 0.)
I_UG15 ( 17 119 ) COMPLEX( 7.53066K, 0.)
I_UG16 ( 14 118 ) COMPLEX( 7.53066K, 0.)
I_UG17 ( 20 128 ) COMPLEX( 7.53066K, 0.)
I_UG18 ( 19 127 ) COMPLEX( 7.53066K, 0.)
I_UG19 ( 21 125 ) COMPLEX( 7.53066K, 0.)
I_UG20 ( 18 124 ) COMPLEX( 7.53066K, 0.)
I_UG21 ( 24 134 ) COMPLEX( 0.3623188, 0.)
I_UG22 ( 23 133 ) COMPLEX( 0.3623188, 0.)
I_UG23 ( 25 131 ) COMPLEX( 0.3623188, 0.)
I_UG24 ( 22 130 ) COMPLEX( 0.3623188, 0.)
I_UG25 ( 28 140 ) COMPLEX( 0.3623188, 0.)
I_UG26 ( 27 139 ) COMPLEX( 0.3623188, 0.)
I_UG27 ( 29 137 ) COMPLEX( 0.3623188, 0.)
I_UG28 ( 26 136 ) COMPLEX( 0.3623188, 0.)
I_UG29 ( 32 158 ) COMPLEX( 0.3623188, 0.)
I_UG30 ( 31 157 ) COMPLEX( 0.3623188, 0.)
I_UG31 ( 33 155 ) COMPLEX( 0.3623188, 0.)
I_UG32 ( 30 154 ) COMPLEX( 0.3623188, 0.)
I_UG33 ( 36 152 ) COMPLEX( 0.3623188, 0.)
I_UG34 ( 35 151 ) COMPLEX( 0.3623188, 0.)
I_UG35 ( 37 149 ) COMPLEX( 0.3623188, 0.)
I_UG36 ( 34 148 ) COMPLEX( 0.3623188, 0.)
I_UG37 ( 40 146 ) COMPLEX( 0.3623188, 0.)
I_UG38 ( 39 145 ) COMPLEX( 0.3623188, 0.)
I_UG39 ( 41 143 ) COMPLEX( 0.3623188, 0.)
I_UG40 ( 38 142 ) COMPLEX( 0.3623188, 0.)
I_UG41 ( 44 98 ) COMPLEX( 7.53066K, 0.)
I_UG42 ( 43 97 ) COMPLEX( 7.53066K, 0.)
I_UG43 ( 45 95 ) COMPLEX( 7.53066K, 0.)
I_UG44 ( 42 94 ) COMPLEX( 7.53066K, 0.)
I_UG45 ( 48 92 ) COMPLEX( 7.53066K, 0.)
I_UG46 ( 47 91 ) COMPLEX( 7.53066K, 0.)
I_UG47 ( 49 89 ) COMPLEX( 7.53066K, 0.)
I_UG48 ( 46 88 ) COMPLEX( 7.53066K, 0.)
I_UG49 ( 161 86 ) COMPLEX( 7.53066K, 0.)
I_UG50 ( 1 84 ) COMPLEX( 7.53066K, 0.)
**** 
* For radial impedance load: 
V_UG05 ( 4 104 ) COMPLEX( 11.8K, 0.) 
V_UG06 ( 3 103 ) COMPLEX( 13.8K, 0.) 
V_UG07 ( 5 101 ) COMPLEX( 13.8K, 0.) 
V_UG08 ( 2 100 ) COMPLEX( 13.8K, 0.) 
V_UG09 ( 12 116 ) COMPLEX( 13.8K, 0.) 
V_UG10 ( 11 115 ) COMPLEX( 13.8K, 0.) 
V_UG11 ( 13 113 ) COMPLEX( 13.8K, 0.) 
V_UG12 ( 10 112 ) COMPLEX( 13.8K, 0.) 
V_UG13 ( 16 122 ) COMPLEX( 13.8K, 0.) 
V_UG14 ( 15 121 ) COMPLEX( 13.8K, 0.) 
V_UG15 ( 17 119 ) COMPLEX( 13.8K, 0.) 
V_UG16 ( 14 118 ) COMPLEX( 13.8K, 0.) 
V_UG17 ( 20 128 ) COMPLEX( 13.8K, 0.) 
V_UG18 ( 19 127 ) COMPLEX( 13.8K, 0.) 
V_UG19 ( 21 125 ) COMPLEX( 13.8K, 0.) 
V_UG20 ( 18 124 ) COMPLEX( 13.8K, 0.) 
V_UG21 ( 24 134 ) COMPLEX( 13.8K, 0.) 
V_UG22 ( 23 133 ) COMPLEX( 13.8K, 0.) 
V_UG23 ( 25 131 ) COMPLEX( 13.8K, 0.) 
V_UG24 ( 22 130 ) COMPLEX( 13.8K, 0.) 
V_UG25 ( 28 140 ) COMPLEX( 13.8K, 0.) 
V_UG26 ( 27 139 ) COMPLEX( 13.8K, 0.) 
V_UG27 ( 29 137 ) COMPLEX( 13.8K, 0.) 
V_UG28 ( 26 136 ) COMPLEX( 13.8K, 0.) 
V_UG29 ( 32 158 ) COMPLEX( 13.8K, 0.) 
V_UG30 ( 31 157 ) COMPLEX( 13.8K, 0.) 
V_UG31 ( 33 155 ) COMPLEX( 13.8K, 0.) 
V_UG32 ( 30 154 ) COMPLEX( 13.8K, 0.) 
V_UG33 ( 36 152 ) COMPLEX( 13.8K, 0.) 
V_UG34 ( 35 151 ) COMPLEX( 13.8K, 0.) 
V_UG35 ( 37 149 ) COMPLEX( 13.8K, 0.) 
V_UG36 ( 34 148 ) COMPLEX( 13.8K, 0.) 
V_UG37 ( 40 146 ) COMPLEX( 13.8K, 0.) 
V_UG38 ( 39 145 ) COMPLEX( 13.8K, 0.) 
V_UG39 ( 41 143 ) COMPLEX( 13.8K, 0.) 
V_UG40 ( 38 142 ) COMPLEX( 13.8K, 0.) 
V_UG41 ( 44 98 ) COMPLEX( 13.8K, 0.) 
V_UG42 ( 43 97 ) COMPLEX( 13.8K, 0.) 
V_UG43 ( 45 95 ) COMPLEX( 13.8K, 0.) 
V_UG44 ( 42 94 ) COMPLEX( 13.8K, 0.) 
V_UG45 ( 48 92 ) COMPLEX( 13.8K, 0.) 
V_UG46 ( 47 91 ) COMPLEX( 13.8K, 0.) 
V_UG47 ( 49 89 ) COMPLEX( 13.8K, 0.) 
V_UG48 ( 46 88 ) COMPLEX( 13.8K, 0.) 
********* Inverted phase (180.0) V_UG49 ( 161 86 ) ( 161 86 ) COMPLEX( 13.8K, 0.) 
*****V_UG49 ( 86 161 ) COMPLEX( 13.8K, 0.) 
********* Inverted phase (180.0) V_UG50 ( 1 84 ) ( 1 84 ) COMPLEX( 13.8K, 0.) 
*****V_UG50 ( 84 1 ) COMPLEX( 13.8K, 0.) 
X_T01 ( 105 108 242 )  MONOPHASIC_TRANSFORMER_525K
X_T02 ( 99 102 244 )  MONOPHASIC_TRANSFORMER_525K
X_T03 ( 111 114 266 )  MONOPHASIC_TRANSFORMER_525K
X_T04 ( 117 120 265 )  MONOPHASIC_TRANSFORMER_525K
X_T05 ( 123 126 263 )  MONOPHASIC_TRANSFORMER_525K
X_T06 ( 129 132 260 )  MONOPHASIC_TRANSFORMER_525K
X_T07 ( 135 138 259 )  MONOPHASIC_TRANSFORMER_525K
X_T08 ( 153 156 257 )  MONOPHASIC_TRANSFORMER_525K
X_T09 ( 147 150 255 )  MONOPHASIC_TRANSFORMER_525K
X_T10 ( 141 144 253 )  MONOPHASIC_TRANSFORMER_525K
X_T11 ( 93 96 250 )  MONOPHASIC_TRANSFORMER_525K
X_T12 ( 87 90 249 )  MONOPHASIC_TRANSFORMER_525K
X_T13 ( 83 85 247 )  MONOPHASIC_TRANSFORMER_525K
***R_LT3_METER ( 52 268 ) COMPLEX( 200.n , 0.) 
***R_LT2_METER ( 54 270 ) COMPLEX( 200.n , 0.) 
R_LT3_METER ( 268 3600 ) COMPLEX( 200.n, 0.)
R_LT3_METER1 ( 52 3599 ) COMPLEX( 100.n, 0.)
R_LT2_METER ( 270 3598 ) COMPLEX( 200.n, 0.)
R_LT2_METER1 ( 54 3597 ) COMPLEX( 100.n, 0.)
R_LT1_METER ( 269 3595 ) COMPLEX( 200.n, 0.)
R_LT1_METER1 ( 53 3596 ) COMPLEX( 100.n, 0.)
* 
X_LT1 ( 3596 3595 )  LT_LT1_LT2
X_LT2 ( 3597 3598 )  LT_LT1_LT2
X_LT3 ( 3599 3600 )  LT_LT3
* 
* Infinite grid/bar; power or current depend on V_Grid: 
**** TEST R_Grid_SWITCH ( 50 273 ) COMPLEX( 100.n, 0.)
R_Grid_SWITCH ( 50 271 ) COMPLEX( 100.n, 0.)
V_Grid ( 271 0 ) COMPLEX( 676.107K,-3.85972K)
* Reactance Xss at the secondary: Xss = 0.43*(525/13.8)^2 = 622.34168241966 
**** TEST R_Grid ( 271 273 ) COMPLEX( 0.0144731, 622.342)
R_Grid ( 0 0 ) COMPLEX( 0.0144731, 622.342)
* 
* Radial. finite grid/bar: 
R_LOAD_BARRA_B ( 0 272 ) COMPLEX( 30.4697K,-217.775)
R_LOAD_BARRA_B_SWITCH ( 0 0 ) COMPLEX( 1.E+12, 0.)
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA Geral 
R_S891xxQCE11 ( 274 368 ) COMPLEX( 100.n, 0.)
R_S891xxQCE12 ( 275 375 ) COMPLEX( 100.n, 0.)
R_D52CARGAxxQCMAC2 ( 0 353 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxQCMAC1 ( 0 525 ) COMPLEX( 387.2, 0.)
****R_D52CARGAxxTSVT2 ( 0 320 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxCDTSB4 ( 0 276 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxTSVT1 ( 0 342 ) COMPLEX( 387.2, 0.)
R_D52CARGAxxCDTSB3 ( 0 277 ) COMPLEX( 387.2, 0.)
****R_D52CARGAxxQCME2 ( 0 432 ) COMPLEX( 387.2, 0.)
R_D52QLxxQCM11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSE3 ( 516 511 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSB2 ( 456 529 )  MONOPHASIC_REGULATOR
X_TSE2 ( 522 526 )  MONOPHASIC_TRANSFORMER_440
R_D52QEExxQCM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE1xxQCM2 ( 531 455 ) COMPLEX( 100.n, 0.)
X_TSA3 ( 530 531 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE2xxQCM2 ( 532 453 ) COMPLEX( 100.n, 0.)
X_TSA4 ( 528 532 )  MONOPHASIC_TRANSFORMER_440
R_D52QLxxQCM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxQCGE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxQCGE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxCDG26 ( 83 387 ) COMPLEX( 100.n, 0.)
R_D52xxCDG25 ( 85 386 ) COMPLEX( 100.n, 0.)
X_TSA26 ( 387 388 )  MONOPHASIC_TRANSFORMER_440
X_TSA25 ( 386 385 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM13 ( 388 389 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM13 ( 385 390 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QLxxQCM13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSE13 ( 383 384 )  MONOPHASIC_TRANSFORMER_440
R_S891xxQCE13 ( 382 383 ) COMPLEX( 100.n, 0.)
R_S892xxQCE13 ( 374 382 ) COMPLEX( 100.n, 0.)
R_S893xxQCE13 ( 381 382 ) COMPLEX( 100.n, 0.)
R_D52206xxQCM13 ( 389 402 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM13 ( 389 406 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM13 ( 395 389 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM13 ( 389 403 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM13 ( 389 404 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM13 ( 405 389 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM13 ( 390 401 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM13 ( 390 399 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM13 ( 390 397 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM13 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQCM13 ( 390 400 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM13 ( 396 390 ) COMPLEX( 100.n, 0.)
R_D52QLxxQCM12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSE7 ( 335 327 )  MONOPHASIC_TRANSFORMER_440
X_TSB4 ( 322 323 )  MONOPHASIC_REGULATOR
R_D52xxCDTSB4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxCDG14E ( 135 324 ) COMPLEX( 100.n, 0.)
R_D522xxCDG14S ( 323 324 ) COMPLEX( 100.n, 0.)
R_D521xxCDG14S ( 324 325 ) COMPLEX( 100.n, 0.)
R_D52xxCDG13 ( 138 326 ) COMPLEX( 100.n, 0.)
R_D52QLxxQCM7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSA14 ( 325 328 )  MONOPHASIC_TRANSFORMER_440
X_TSA13 ( 326 329 )  MONOPHASIC_TRANSFORMER_440
X_TSVT2 ( 320 321 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM7 ( 328 330 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM7 ( 329 331 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQCM7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQCM7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQCM7 ( 330 554 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM7 ( 552 330 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM7 ( 330 553 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM7 ( 330 551 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM7 ( 331 550 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM7 ( 331 548 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM7 ( 331 546 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM7 ( 547 331 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM7 ( 331 549 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207xxQCM6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSVT1 ( 342 341 )  MONOPHASIC_TRANSFORMER_440
X_TSE6 ( 337 338 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDTSB3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSB3 ( 348 349 )  MONOPHASIC_REGULATOR
R_D522xxCDG12S ( 347 348 ) COMPLEX( 100.n, 0.)
R_D521xxCDG12S ( 346 347 ) COMPLEX( 100.n, 0.)
R_D52ExxCDG12E ( 129 347 ) COMPLEX( 100.n, 0.)
X_TSA12 ( 346 345 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM6 ( 345 343 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM6 ( 340 344 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QLxxQCM6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSA11 ( 339 340 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG11 ( 132 339 ) COMPLEX( 100.n, 0.)
R_D52206xxQCM6 ( 343 555 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQCM6 ( 343 566 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM6 ( 564 343 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM6 ( 343 565 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM6 ( 343 562 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM6 ( 344 561 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM6 ( 344 559 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM6 ( 344 557 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM6 ( 558 344 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM6 ( 344 560 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQCM5 ( 449 567 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM5 ( 449 578 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM5 ( 449 574 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQCM5 ( 576 449 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM5 ( 449 577 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM5 ( 450 573 ) COMPLEX( 100.n, 0.)
R_D52QLxxQCM5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQCM5 ( 450 571 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM5 ( 450 569 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM5 ( 570 450 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM5 ( 450 572 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSE5 ( 333 315 )  MONOPHASIC_TRANSFORMER_440
* X_TSG1 ( 351 437 ) MONOPHASIC_TRANSFORMER_440 
X_TSG1 ( 437 351 )  MONOPHASIC_TRANSFORMER_440
X_TSG2 ( 436 350 )  MONOPHASIC_TRANSFORMER_440
R_S892xxQCE11 ( 366 274 ) COMPLEX( 100.n, 0.)
R_S893xxQCE11 ( 274 367 ) COMPLEX( 100.n, 0.)
X_TSE11 ( 368 369 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM11 ( 373 364 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE1xxQCM11 ( 370 365 ) COMPLEX( 100.n, 0.)
X_TSA21 ( 371 370 )  MONOPHASIC_TRANSFORMER_440
X_TSA22 ( 372 373 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG21 ( 96 371 ) COMPLEX( 100.n, 0.)
R_D52xxCDG22 ( 93 372 ) COMPLEX( 100.n, 0.)
V_UGD7 ( 391 0 ) COMPLEX( 255.7662, 0.)
R_UGD7 ( 3728 3720 ) COMPLEX( 100.n, 0.)
R_D52xxQCGE7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSG7 ( 393 392 )  MONOPHASIC_TRANSFORMER_440
R_D522xxQCME4 ( 393 394 ) COMPLEX( 100.n, 0.)
R_D523xxQCME4 ( 394 381 ) COMPLEX( 100.n, 0.)
R_D521xxQCME4 ( 394 439 ) COMPLEX( 100.n, 0.)
R_D52QLxxQCM3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QEExxQCM3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE1xxQCM3 ( 513 425 ) COMPLEX( 100.n, 0.)
X_TSA5 ( 521 513 )  MONOPHASIC_TRANSFORMER_440
X_TSA6 ( 514 512 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM3 ( 512 424 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE1xxQCM4 ( 506 452 ) COMPLEX( 100.n, 0.)
X_TSE4 ( 509 504 )  MONOPHASIC_TRANSFORMER_440
X_TSA7 ( 510 506 )  MONOPHASIC_TRANSFORMER_440
X_TSB6 ( 441 459 )  MONOPHASIC_REGULATOR
R_D52QLxxQCM10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QLxxQCM9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QLxxQCM4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE2xxQCM4 ( 505 451 ) COMPLEX( 100.n, 0.)
X_TSA8 ( 507 505 )  MONOPHASIC_TRANSFORMER_440
R_S891xxQCE8 ( 502 503 ) COMPLEX( 100.n, 0.)
R_S892xxQCE8 ( 440 502 ) COMPLEX( 100.n, 0.)
R_S893xxQCE8 ( 442 502 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM11 ( 365 538 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM11 ( 365 534 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM11 ( 365 536 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM11 ( 364 539 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM11 ( 542 364 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM11 ( 364 541 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM11 ( 364 540 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM11 ( 364 543 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM11 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQCM11 ( 365 537 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM11 ( 533 365 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM12 ( 363 413 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM12 ( 363 409 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM12 ( 363 411 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM12 ( 362 414 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM12 ( 417 362 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM12 ( 362 416 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM12 ( 362 415 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM12 ( 362 418 ) COMPLEX( 100.n, 0.)
R_D52206xxQCM12 ( 407 362 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQCM12 ( 363 412 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM12 ( 408 363 ) COMPLEX( 100.n, 0.)
R_S893xxQCE12 ( 275 374 ) COMPLEX( 100.n, 0.)
R_S892xxQCE12 ( 367 275 ) COMPLEX( 100.n, 0.)
X_TSE12 ( 375 376 )  MONOPHASIC_TRANSFORMER_440
R_D52QEExxQCM12 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE1xxQCM12 ( 377 363 ) COMPLEX( 100.n, 0.)
R_D52QE2xxQCM12 ( 380 362 ) COMPLEX( 100.n, 0.)
X_TSA24 ( 379 380 )  MONOPHASIC_TRANSFORMER_440
X_TSA23 ( 378 377 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG24 ( 87 379 ) COMPLEX( 100.n, 0.)
R_D52xxCDG23 ( 90 378 ) COMPLEX( 100.n, 0.)
V_UGD5 ( 355 0 ) COMPLEX( 255.7662, 0.)
*RUGD5n ( 355 3726 ) FIT (1,1 227.73,5 281.082645,210 338.264463,430) order = 1
R_UGD5 ( 3726 3718 ) COMPLEX( 100.n, 0.)
V_UGD6 ( 356 0 ) COMPLEX( 255.7662, 0.)
*RUGD6n ( 356 3727 ) FIT (1,1 227.73,5 281.082645,210 338.264463,430) order = 1
R_UGD6 ( 3727 3719 ) COMPLEX( 100.n, 0.)
R_D52xxQCGE5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxQCGE6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSG5 ( 360 357 )  MONOPHASIC_TRANSFORMER_440
X_TSG6 ( 359 358 )  MONOPHASIC_TRANSFORMER_440
R_D525xxQCME3 ( 361 439 ) COMPLEX( 100.n, 0.)
R_D522xxQCME3 ( 361 440 ) COMPLEX( 100.n, 0.)
R_D524xxQCME3 ( 359 361 ) COMPLEX( 100.n, 0.)
R_D523xxQCME3 ( 360 361 ) COMPLEX( 100.n, 0.)
R_D521xxQCME3 ( 354 361 ) COMPLEX( 100.n, 0.)
R_D525Q1xxQCMAC2 ( 353 441 ) COMPLEX( 100.n, 0.)
R_D524Q1xxQCMAC2 ( 353 354 ) COMPLEX( 100.n, 0.)
R_D522Q1xxQCMAC2 ( 354 445 ) COMPLEX( 100.n, 0.)
R_D525xxQCME2 ( 307 435 ) COMPLEX( 100.n, 0.)
R_D521xxQCME2 ( 435 427 ) COMPLEX( 100.n, 0.)
R_D524xxQCME2 ( 432 435 ) COMPLEX( 100.n, 0.)
R_D523xxQCME2 ( 433 435 ) COMPLEX( 100.n, 0.)
R_D522xxQCME2 ( 434 435 ) COMPLEX( 100.n, 0.)
X_TSG3 ( 434 430 )  MONOPHASIC_TRANSFORMER_440
X_TSG4 ( 433 431 )  MONOPHASIC_TRANSFORMER_440
R_D52xxQCGE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxQCGE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
V_UGD4 ( 428 0 ) COMPLEX( 255.7662, 0.)
R_UGD4 ( 3725 3717 ) COMPLEX( 100.n, 0.)
V_UGD3 ( 429 0 ) COMPLEX( 255.7662, 0.)
R_UGD3 ( 3724 3716 ) COMPLEX( 100.n, 0.)
V_UGD2 ( 352 0 ) COMPLEX( 255.7662, 0.)
R_UGD2 ( 3723 3715 ) COMPLEX( 100.n, 0.)
V_UGD1 ( 527 0 ) COMPLEX( 255.7662, 0.)
R_UGD1 ( 3722 3714 ) COMPLEX( 100.n, 0.)
R_D524xxQCME1 ( 436 438 ) COMPLEX( 100.n, 0.)
R_D523xxQCME1 ( 437 438 ) COMPLEX( 100.n, 0.)
R_D525xxQCME1 ( 427 438 ) COMPLEX( 100.n, 0.)
R_D522xxQCME1 ( 438 313 ) COMPLEX( 100.n, 0.)
R_D521xxQCME1 ( 314 438 ) COMPLEX( 100.n, 0.)
R_D524Q1xxQCMAC1 ( 314 525 ) COMPLEX( 100.n, 0.)
R_D525Q1xxQCMAC1 ( 525 456 ) COMPLEX( 100.n, 0.)
R_D522Q1xxQCMAC1 ( 524 314 ) COMPLEX( 100.n, 0.)
R_D52ExxCDG20E ( 141 460 ) COMPLEX( 100.n, 0.)
R_D522xxCDG20S ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D521xxCDG20S ( 460 461 ) COMPLEX( 100.n, 0.)
R_D52xxCDG19 ( 144 467 ) COMPLEX( 100.n, 0.)
X_TSA20 ( 461 463 )  MONOPHASIC_TRANSFORMER_440
X_TSA19 ( 467 464 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM10 ( 463 419 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM10 ( 464 420 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQCM10 ( 419 458 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM10 ( 419 482 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM10 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQCM10 ( 419 483 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM10 ( 484 419 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM10 ( 419 481 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM10 ( 420 480 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM10 ( 420 478 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM10 ( 420 476 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM10 ( 477 420 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM10 ( 420 479 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM10 ( 475 420 ) COMPLEX( 100.n, 0.)
R_D52xxCDG18 ( 147 471 ) COMPLEX( 100.n, 0.)
R_D52xxCDG17 ( 150 474 ) COMPLEX( 100.n, 0.)
R_S892xxQCE9 ( 442 472 ) COMPLEX( 100.n, 0.)
R_S893xxQCE9 ( 457 472 ) COMPLEX( 100.n, 0.)
R_S891xxQCE9 ( 472 473 ) COMPLEX( 100.n, 0.)
R_S892xxQCE10 ( 457 465 ) COMPLEX( 100.n, 0.)
R_S893xxQCE10 ( 366 465 ) COMPLEX( 100.n, 0.)
R_S891xxQCE10 ( 465 466 ) COMPLEX( 100.n, 0.)
X_TSE10 ( 466 462 )  MONOPHASIC_TRANSFORMER_440
X_TSE9 ( 473 468 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM9 ( 469 422 ) COMPLEX( 100.n, 0.)
X_TSA18 ( 471 469 )  MONOPHASIC_TRANSFORMER_440
X_TSA17 ( 474 470 )  MONOPHASIC_TRANSFORMER_440
R_D52QE1xxQCM9 ( 470 423 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM9 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQCM9 ( 421 422 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM9 ( 422 493 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM9 ( 422 496 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM9 ( 422 494 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM9 ( 495 422 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM9 ( 422 492 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM9 ( 423 491 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM9 ( 423 489 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM9 ( 423 487 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM9 ( 488 423 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM9 ( 423 490 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM9 ( 486 423 ) COMPLEX( 100.n, 0.)
X_TSB5 ( 445 447 )  MONOPHASIC_REGULATOR
X_TSE8 ( 503 497 )  MONOPHASIC_TRANSFORMER_440
R_D52QE2xxQCM8 ( 498 443 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM8 ( 499 444 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM8 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSA16 ( 500 498 )  MONOPHASIC_TRANSFORMER_440
X_TSA15 ( 448 499 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG16 ( 153 500 ) COMPLEX( 100.n, 0.)
R_D522xxCDG15S ( 446 448 ) COMPLEX( 100.n, 0.)
R_D521xxCDG15S ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxCDG15E ( 156 446 ) COMPLEX( 100.n, 0.)
R_D52xxCDG8 ( 117 507 ) COMPLEX( 100.n, 0.)
R_D52xxCDG7 ( 120 510 ) COMPLEX( 100.n, 0.)
R_D52xxCDG6 ( 111 514 ) COMPLEX( 100.n, 0.)
R_D52xxCDG5 ( 114 521 ) COMPLEX( 100.n, 0.)
R_D52206xxQCM2 ( 454 453 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQCM2 ( 453 589 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM2 ( 587 453 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM2 ( 453 588 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM2 ( 453 585 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM2 ( 455 584 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM2 ( 455 582 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM2 ( 455 580 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM2 ( 581 455 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM2 ( 455 583 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM2 ( 579 455 ) COMPLEX( 100.n, 0.)
R_D52QE2xxQCM5 ( 318 449 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM5 ( 319 450 ) COMPLEX( 100.n, 0.)
R_D52QEExxQCM5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSA10 ( 317 318 )  MONOPHASIC_TRANSFORMER_440
X_TSA9 ( 316 319 )  MONOPHASIC_TRANSFORMER_440
R_D52xxCDG10 ( 123 317 ) COMPLEX( 100.n, 0.)
R_D52xxCDG9 ( 126 316 ) COMPLEX( 100.n, 0.)
R_S893xxQCE6 ( 306 336 ) COMPLEX( 100.n, 0.)
R_C574xxQCE6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE6 ( 308 336 ) COMPLEX( 100.n, 0.)
R_C573xxQCE6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE6 ( 336 337 ) COMPLEX( 100.n, 0.)
R_C571xxQCE6 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE7 ( 306 334 ) COMPLEX( 100.n, 0.)
R_C574xxQCE7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE7 ( 307 334 ) COMPLEX( 100.n, 0.)
R_C573xxQCE7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE7 ( 334 335 ) COMPLEX( 100.n, 0.)
R_C571xxQCE7 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE5 ( 308 332 ) COMPLEX( 100.n, 0.)
R_C574xxQCE5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE5 ( 309 332 ) COMPLEX( 100.n, 0.)
R_C573xxQCE5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE5 ( 332 333 ) COMPLEX( 100.n, 0.)
R_C571xxQCE5 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE2 ( 311 520 ) COMPLEX( 100.n, 0.)
R_C574xxQCE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE2 ( 312 520 ) COMPLEX( 100.n, 0.)
R_C573xxQCE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE2 ( 520 522 ) COMPLEX( 100.n, 0.)
R_C571xxQCE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE3 ( 310 515 ) COMPLEX( 100.n, 0.)
R_C574xxQCE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE3 ( 311 515 ) COMPLEX( 100.n, 0.)
R_C573xxQCE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE3 ( 515 516 ) COMPLEX( 100.n, 0.)
R_C571xxQCE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE4 ( 309 508 ) COMPLEX( 100.n, 0.)
R_C574xxQCE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE4 ( 310 508 ) COMPLEX( 100.n, 0.)
R_C573xxQCE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE4 ( 508 509 ) COMPLEX( 100.n, 0.)
R_C571xxQCE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S893xxQCE1 ( 312 517 ) COMPLEX( 100.n, 0.)
R_C574xxQCE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S892xxQCE1 ( 313 517 ) COMPLEX( 100.n, 0.)
R_C573xxQCE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_C572xxQCE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_S891xxQCE1 ( 517 518 ) COMPLEX( 100.n, 0.)
R_C571xxQCE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
X_TSE1 ( 518 519 )  MONOPHASIC_TRANSFORMER_440
R_D52201xxQCM3 ( 424 597 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM3 ( 424 601 ) COMPLEX( 100.n, 0.)
R_D52206xxQCM3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQCM3 ( 424 598 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM3 ( 599 424 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM3 ( 424 600 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM3 ( 425 596 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM3 ( 425 594 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM3 ( 425 592 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM3 ( 593 425 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM3 ( 425 595 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQCM4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQCM4 ( 451 622 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM4 ( 620 451 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM4 ( 451 621 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM4 ( 451 618 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM4 ( 452 616 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM4 ( 452 614 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM4 ( 615 452 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM4 ( 452 617 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQCM8 ( 443 609 ) COMPLEX( 100.n, 0.)
R_D52205xxQCM8 ( 443 612 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM8 ( 443 610 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM8 ( 611 443 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM8 ( 443 608 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM8 ( 444 607 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM8 ( 444 605 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM8 ( 444 603 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM8 ( 604 444 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM8 ( 444 606 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM8 ( 602 444 ) COMPLEX( 100.n, 0.)
R_D52204xxQCM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQCM1 ( 624 638 ) COMPLEX( 100.n, 0.)
R_D52203xxQCM1 ( 624 636 ) COMPLEX( 100.n, 0.)
R_D52202xxQCM1 ( 637 624 ) COMPLEX( 100.n, 0.)
R_D52201xxQCM1 ( 624 634 ) COMPLEX( 100.n, 0.)
R_D52106xxQCM1 ( 623 633 ) COMPLEX( 100.n, 0.)
R_D52105xxQCM1 ( 623 630 ) COMPLEX( 100.n, 0.)
R_D52104xxQCM1 ( 623 626 ) COMPLEX( 100.n, 0.)
R_D52103xxQCM1 ( 629 623 ) COMPLEX( 100.n, 0.)
R_D52102xxQCM1 ( 623 632 ) COMPLEX( 100.n, 0.)
R_D52101xxQCM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QEExxQCM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52QE2xxQCM1 ( 631 624 ) COMPLEX( 100.n, 0.)
R_D52QE1xxQCM1 ( 628 623 ) COMPLEX( 100.n, 0.)
X_TSA2 ( 627 631 )  MONOPHASIC_TRANSFORMER_440
X_TSA1 ( 523 628 )  MONOPHASIC_TRANSFORMER_440
X_TSB1 ( 426 524 )  MONOPHASIC_REGULATOR
R_D52ExxCDG3E ( 102 302 ) COMPLEX( 100.n, 0.)
R_D522xxCDG3S ( 302 530 ) COMPLEX( 100.n, 0.)
R_D521xxCDG3S ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52xxCDG4 ( 99 528 ) COMPLEX( 100.n, 0.)
R_D52xxCDG2 ( 105 627 ) COMPLEX( 100.n, 0.)
R_D521xxCDG1S ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D522xxCDG1S ( 303 523 ) COMPLEX( 100.n, 0.)
R_D52ExxCDG1E ( 108 303 ) COMPLEX( 100.n, 0.)
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG1 
R_D52322LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52322xxQSG1 ( 639 640 ) COMPLEX( 100.n, 0.)
R_D52323LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52323xxQSG1 ( 641 640 ) COMPLEX( 100.n, 0.)
R_D52321LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52321xxQSG1 ( 642 640 ) COMPLEX( 100.n, 0.)
R_D52320LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52320xxQSG1 ( 640 643 ) COMPLEX( 100.n, 0.)
R_D52307xxQSG1 ( 644 640 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309xxQSG1 ( 645 640 ) COMPLEX( 100.n, 0.)
R_D52309LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319xxQSG1 ( 646 640 ) COMPLEX( 100.n, 0.)
R_D52318LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52318xxQSG1 ( 647 640 ) COMPLEX( 100.n, 0.)
R_D52310LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52310xxQSG1 ( 648 640 ) COMPLEX( 100.n, 0.)
R_D52317LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52317xxQSG1 ( 649 640 ) COMPLEX( 100.n, 0.)
R_D52316LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52316xxQSG1 ( 650 640 ) COMPLEX( 100.n, 0.)
R_D52315LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52315xxQSG1 ( 651 640 ) COMPLEX( 100.n, 0.)
R_D52314LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52314xxQSG1 ( 652 640 ) COMPLEX( 100.n, 0.)
R_D52313LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52313xxQSG1 ( 653 640 ) COMPLEX( 100.n, 0.)
R_D52312LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52312xxQSG1 ( 654 640 ) COMPLEX( 100.n, 0.)
R_D52311LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52311xxQSG1 ( 655 640 ) COMPLEX( 100.n, 0.)
R_D52308xxQSG1 ( 656 640 ) COMPLEX( 100.n, 0.)
R_D52308LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSG1 ( 657 640 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSG1 ( 658 640 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSG1 ( 659 640 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSG1 ( 660 640 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSG1 ( 661 640 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSG1 ( 640 662 ) COMPLEX( 100.n, 0.)
R_D52207xxQSG1 ( 664 665 ) COMPLEX( 100.n, 0.)
R_D52207LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52209xxQSG1 ( 666 665 ) COMPLEX( 100.n, 0.)
R_D52209LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52219LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52219xxQSG1 ( 667 665 ) COMPLEX( 100.n, 0.)
R_D52218LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52218xxQSG1 ( 668 665 ) COMPLEX( 100.n, 0.)
R_D52210LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52210xxQSG1 ( 669 665 ) COMPLEX( 100.n, 0.)
R_D52217LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52217xxQSG1 ( 670 665 ) COMPLEX( 100.n, 0.)
R_D52216LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52216xxQSG1 ( 671 665 ) COMPLEX( 100.n, 0.)
R_D52215LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52215xxQSG1 ( 672 665 ) COMPLEX( 100.n, 0.)
R_D52214LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52214xxQSG1 ( 673 665 ) COMPLEX( 100.n, 0.)
R_D52213LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52213xxQSG1 ( 674 665 ) COMPLEX( 100.n, 0.)
R_D52212LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52212xxQSG1 ( 675 665 ) COMPLEX( 100.n, 0.)
R_D52211LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52211xxQSG1 ( 676 665 ) COMPLEX( 100.n, 0.)
R_D52208xxQSG1 ( 677 665 ) COMPLEX( 100.n, 0.)
R_D52208LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQSG1 ( 678 665 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQSG1 ( 679 665 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQSG1 ( 680 665 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSG1 ( 681 665 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSG1 ( 682 665 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSG1 ( 665 683 ) COMPLEX( 100.n, 0.)
R_D52E1xxQSG1 ( 626 687 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSG1 ( 585 665 ) COMPLEX( 100.n, 0.)
R_D52L2xxQSG1 ( 640 665 ) COMPLEX( 100.n, 0.)
R_D52107xxQSG1 ( 686 687 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSG1 ( 688 687 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxQSG1 ( 689 687 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxQSG1 ( 690 687 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxQSG1 ( 691 687 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxQSG1 ( 692 687 ) COMPLEX( 100.n, 0.)
R_D52L1xxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxQSG1 ( 694 687 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSG1 ( 695 687 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxQSG1 ( 696 687 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSG1 ( 697 687 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSG1 ( 698 687 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxQSG1 ( 699 687 ) COMPLEX( 100.n, 0.)
R_D52108xxQSG1 ( 700 687 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSG1 ( 701 687 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSG1 ( 702 687 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSG1 ( 703 687 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSG1 ( 704 687 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSG1 ( 705 687 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSG1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSG1 ( 687 706 ) COMPLEX( 100.n, 0.)
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG2 
R_D52207xxQSG2 ( 708 709 ) COMPLEX( 100.n, 0.)
R_D52207LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52209xxQSG2 ( 710 709 ) COMPLEX( 100.n, 0.)
R_D52209LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52210LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52210xxQSG2 ( 711 709 ) COMPLEX( 100.n, 0.)
R_D52216LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52216xxQSG2 ( 712 709 ) COMPLEX( 100.n, 0.)
R_D52215LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52215xxQSG2 ( 713 709 ) COMPLEX( 100.n, 0.)
R_D52214LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52214xxQSG2 ( 714 709 ) COMPLEX( 100.n, 0.)
R_D52213LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52213xxQSG2 ( 715 709 ) COMPLEX( 100.n, 0.)
R_D52212LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52212xxQSG2 ( 716 709 ) COMPLEX( 100.n, 0.)
R_D52211LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52211xxQSG2 ( 717 709 ) COMPLEX( 100.n, 0.)
R_D52208xxQSG2 ( 718 709 ) COMPLEX( 100.n, 0.)
R_D52208LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQSG2 ( 719 709 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQSG2 ( 720 709 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQSG2 ( 721 709 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSG2 ( 722 709 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSG2 ( 723 709 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSG2 ( 709 724 ) COMPLEX( 100.n, 0.)
R_D52307xxQSG2 ( 725 726 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309xxQSG2 ( 727 726 ) COMPLEX( 100.n, 0.)
R_D52309LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319xxQSG2 ( 728 726 ) COMPLEX( 100.n, 0.)
R_D52318LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52318xxQSG2 ( 729 726 ) COMPLEX( 100.n, 0.)
R_D52310LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52310xxQSG2 ( 730 726 ) COMPLEX( 100.n, 0.)
R_D52317LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52317xxQSG2 ( 731 726 ) COMPLEX( 100.n, 0.)
R_D52316LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52316xxQSG2 ( 732 726 ) COMPLEX( 100.n, 0.)
R_D52315LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52315xxQSG2 ( 733 726 ) COMPLEX( 100.n, 0.)
R_D52314LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52314xxQSG2 ( 734 726 ) COMPLEX( 100.n, 0.)
R_D52313LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52313xxQSG2 ( 735 726 ) COMPLEX( 100.n, 0.)
R_D52312LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52312xxQSG2 ( 736 726 ) COMPLEX( 100.n, 0.)
R_D52311LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52311xxQSG2 ( 737 726 ) COMPLEX( 100.n, 0.)
R_D52308xxQSG2 ( 738 726 ) COMPLEX( 100.n, 0.)
R_D52308LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSG2 ( 739 726 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSG2 ( 740 726 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSG2 ( 741 726 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSG2 ( 742 726 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSG2 ( 743 726 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSG2 ( 726 744 ) COMPLEX( 100.n, 0.)
R_D52E1xxQSG2 ( 580 748 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSG2 ( 634 709 ) COMPLEX( 100.n, 0.)
R_D52L2xxQSG2 ( 726 709 ) COMPLEX( 100.n, 0.)
R_D52107xxQSG2 ( 747 748 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSG2 ( 749 748 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxQSG2 ( 750 748 ) COMPLEX( 100.n, 0.)
R_D52L1xxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxQSG2 ( 752 748 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSG2 ( 753 748 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxQSG2 ( 754 748 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSG2 ( 755 748 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSG2 ( 756 748 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxQSG2 ( 757 748 ) COMPLEX( 100.n, 0.)
R_D52108xxQSG2 ( 758 748 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSG2 ( 759 748 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSG2 ( 760 748 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSG2 ( 761 748 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSG2 ( 762 748 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSG2 ( 763 748 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSG2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSG2 ( 748 764 ) COMPLEX( 100.n, 0.)
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U01CCM 
R_D52132LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU01 ( 765 766 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU01 ( 767 766 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU01 ( 769 766 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU01 ( 770 766 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU01 ( 771 766 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU01 ( 772 766 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU01 ( 773 766 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125xxU01 ( 774 766 ) COMPLEX( 100.n, 0.)
R_D52124xxU01 ( 775 766 ) COMPLEX( 100.n, 0.)
R_D52117xxU01 ( 776 766 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU01 ( 777 766 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU01 ( 778 766 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU01 ( 779 766 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU01 ( 780 766 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU01 ( 781 766 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU01 ( 766 783 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxU01 ( 784 766 ) COMPLEX( 100.n, 0.)
R_D52ExxU01 ( 630 766 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU01 ( 786 766 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU01 ( 787 766 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU01 ( 788 766 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU01 ( 789 766 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU01 ( 790 766 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU01 ( 791 766 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxU01 ( 792 766 ) COMPLEX( 100.n, 0.)
R_D52107xxU01 ( 793 766 ) COMPLEX( 100.n, 0.)
R_D52108xxU01 ( 794 766 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU01 ( 795 766 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU01 ( 796 766 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU01 ( 797 766 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU01 ( 798 766 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU01 ( 799 766 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU01 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxU01 ( 766 800 ) COMPLEX( 100.n, 0.)
* -------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U02CCM 
R_D52132LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU02 ( 803 802 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU02 ( 807 802 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124xxU02 ( 810 802 ) COMPLEX( 100.n, 0.)
R_D52117xxU02 ( 811 802 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU02 ( 814 802 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU02 ( 816 802 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU02 ( 802 817 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxU02 ( 818 802 ) COMPLEX( 100.n, 0.)
R_D52ExxU02 ( 633 802 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU02 ( 821 802 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU02 ( 822 802 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU02 ( 823 802 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU02 ( 825 802 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxU02 ( 827 802 ) COMPLEX( 100.n, 0.)
R_D52108xxU02 ( 828 802 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU02 ( 830 802 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU02 ( 831 802 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101LOADxxU02 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxU02 ( 802 834 ) COMPLEX( 100.n, 0.)
*------------------------------------------------------------------------------------------------------------------------ 
* Netlist: Auxiliares CA U03CCM 
R_D52132LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU03 ( 835 836 ) COMPLEX( 1.E+12, 0.)
R_D52131LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU03 ( 837 836 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU03 ( 838 836 ) COMPLEX( 1.E+12, 0.)
R_D52129LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU03 ( 839 836 ) COMPLEX( 1.E+12, 0.)
R_D52128LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU03 ( 840 836 ) COMPLEX( 1.E+12, 0.)
R_D52127LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU03 ( 841 836 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU03 ( 842 836 ) COMPLEX( 1.E+12, 0.)
R_D52125LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125xxU03 ( 843 836 ) COMPLEX( 1.E+12, 0.)
R_D52124xxU03 ( 844 836 ) COMPLEX( 100.n, 0.)
R_D52117xxU03 ( 845 836 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU03 ( 846 836 ) COMPLEX( 1.E+12, 0.)
R_D52122LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU03 ( 847 836 ) COMPLEX( 1.E+12, 0.)
R_D52121LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU03 ( 848 836 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU03 ( 849 836 ) COMPLEX( 1.E+12, 0.)
R_D52119LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU03 ( 850 836 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU03 ( 836 851 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxU03 ( 852 836 ) COMPLEX( 100.n, 0.)
R_D52ExxU03 ( 637 836 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU03 ( 854 836 ) COMPLEX( 1.E+12, 0.)
R_D52114LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU03 ( 855 836 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU03 ( 856 836 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU03 ( 857 836 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU03 ( 858 836 ) COMPLEX( 1.E+12, 0.)
R_D52110LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU03 ( 859 836 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxU03 ( 860 836 ) COMPLEX( 1.E+12, 0.)
R_D52107xxU03 ( 861 836 ) COMPLEX( 100.n, 0.)
R_D52108xxU03 ( 862 836 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU03 ( 863 836 ) COMPLEX( 1.E+12, 0.)
R_D52105LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU03 ( 864 836 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU03 ( 865 836 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU03 ( 866 836 ) COMPLEX( 1.E+12, 0.)
R_D52102LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU03 ( 867 836 ) COMPLEX( 1.E+12, 0.)
R_D52101LOADxxU03 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxU03 ( 836 868 ) COMPLEX( 100.n, 0.)
*---------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U04CCM 
R_D52101xxU04 ( 870 902 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU04 ( 901 870 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU04 ( 900 870 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU04 ( 899 870 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU04 ( 898 870 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU04 ( 897 870 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxU04 ( 896 870 ) COMPLEX( 100.n, 0.)
R_D52107xxU04 ( 895 870 ) COMPLEX( 100.n, 0.)
R_D52109xxU04 ( 894 870 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU04 ( 893 870 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU04 ( 892 870 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU04 ( 891 870 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU04 ( 890 870 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU04 ( 889 870 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU04 ( 888 870 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxU04 ( 636 870 ) COMPLEX( 100.n, 0.)
R_D52115xxU04 ( 886 870 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU04 ( 870 885 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU04 ( 884 870 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU04 ( 883 870 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU04 ( 882 870 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU04 ( 881 870 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU04 ( 880 870 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxU04 ( 879 870 ) COMPLEX( 100.n, 0.)
R_D52124xxU04 ( 878 870 ) COMPLEX( 100.n, 0.)
R_D52125xxU04 ( 877 870 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU04 ( 876 870 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU04 ( 875 870 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU04 ( 874 870 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU04 ( 873 870 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU04 ( 872 870 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU04 ( 871 870 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU04 ( 869 870 ) COMPLEX( 100.n, 0.)
R_D52132LOADxxU04 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*--------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSSE1 
R_D52E1xxQSSE1 ( 629 905 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSSE1 ( 589 909 ) COMPLEX( 100.n, 0.)
R_D52307xxQSSE1 ( 918 903 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSSE1 ( 917 903 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSSE1 ( 916 903 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSSE1 ( 915 903 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSSE1 ( 914 903 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSSE1 ( 913 903 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSSE1 ( 912 903 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSSE1 ( 911 909 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSSE1 ( 910 909 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSSE1 ( 908 909 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSSE1 ( 907 905 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSSE1 ( 906 905 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSSE1 ( 904 905 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSSE1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L2xxQSSE1 ( 903 909 ) COMPLEX( 100.n, 0.)
*-------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSSE2 
R_D52E1xxQSSE2 ( 581 921 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSSE2 ( 638 925 ) COMPLEX( 100.n, 0.)
R_D52306xxQSSE2 ( 933 919 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSSE2 ( 932 919 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSSE2 ( 931 919 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSSE2 ( 930 919 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSSE2 ( 929 919 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSSE2 ( 928 919 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSSE2 ( 927 925 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSSE2 ( 926 925 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSSE2 ( 924 925 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSSE2 ( 923 921 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSSE2 ( 922 921 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSSE2 ( 920 921 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSSE2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L2xxQSSE2 ( 919 925 ) COMPLEX( 100.n, 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSAM1 
R_D52101xxQSAM1 ( 935 964 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSAM1 ( 963 935 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSAM1 ( 962 935 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSAM1 ( 961 935 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSAM1 ( 960 935 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSAM1 ( 959 935 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxQSAM1 ( 958 935 ) COMPLEX( 100.n, 0.)
R_D52108xxQSAM1 ( 957 935 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSAM1 ( 956 935 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxQSAM1 ( 955 935 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxQSAM1 ( 954 935 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSAM1 ( 953 935 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSAM1 ( 952 935 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxQSAM1 ( 632 935 ) COMPLEX( 100.n, 0.)
R_D52114xxQSAM1 ( 950 935 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxQSAM1 ( 935 949 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxQSAM1 ( 948 935 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxQSAM1 ( 947 935 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxQSAM1 ( 946 935 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxQSAM1 ( 945 935 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxQSAM1 ( 944 935 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSAM1 ( 943 935 ) COMPLEX( 100.n, 0.)
R_D52122xxQSAM1 ( 942 935 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxQSAM1 ( 941 935 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124xxQSAM1 ( 940 935 ) COMPLEX( 100.n, 0.)
R_D52124LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125xxQSAM1 ( 939 935 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxQSAM1 ( 938 935 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxQSAM1 ( 937 935 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxQSAM1 ( 936 935 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxQSAM1 ( 934 935 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxQSAM1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSAM2 
R_D52101xxQSAM2 ( 975 991 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSAM2 ( 990 975 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSAM2 ( 989 975 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSAM2 ( 988 975 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSAM2 ( 987 975 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSAM2 ( 986 975 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxQSAM2 ( 985 975 ) COMPLEX( 100.n, 0.)
R_D52108xxQSAM2 ( 984 975 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSAM2 ( 983 975 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxQSAM2 ( 982 975 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxQSAM2 ( 981 975 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSAM2 ( 980 975 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSAM2 ( 979 975 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxQSAM2 ( 549 975 ) COMPLEX( 100.n, 0.)
R_D52114xxQSAM2 ( 977 975 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxQSAM2 ( 975 976 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxQSAM2 ( 974 975 ) COMPLEX( 100.n, 0.)
R_D52117LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxQSAM2 ( 973 975 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxQSAM2 ( 972 975 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxQSAM2 ( 971 975 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxQSAM2 ( 970 975 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSAM2 ( 969 975 ) COMPLEX( 100.n, 0.)
R_D52122xxQSAM2 ( 968 975 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxQSAM2 ( 967 975 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124xxQSAM2 ( 966 975 ) COMPLEX( 100.n, 0.)
R_D52124LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52125xxQSAM2 ( 965 975 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxQSAM2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U05CCM 
R_D52101xxU05 ( 993 1025 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU05 ( 1024 993 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU05 ( 1023 993 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU05 ( 1022 993 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU05 ( 1021 993 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU05 ( 1020 993 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxU05 ( 1019 993 ) COMPLEX( 100.n, 0.)
R_D52107xxU05 ( 1018 993 ) COMPLEX( 100.n, 0.)
R_D52109xxU05 ( 1017 993 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU05 ( 1016 993 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU05 ( 1015 993 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU05 ( 1014 993 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU05 ( 1013 993 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU05 ( 1012 993 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU05 ( 1011 993 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxU05 ( 582 993 ) COMPLEX( 100.n, 0.)
R_D52115xxU05 ( 1009 993 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU05 ( 993 1008 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU05 ( 1007 993 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU05 ( 1006 993 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU05 ( 1005 993 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU05 ( 1004 993 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU05 ( 1003 993 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxU05 ( 1002 993 ) COMPLEX( 100.n, 0.)
R_D52124xxU05 ( 1001 993 ) COMPLEX( 100.n, 0.)
R_D52125xxU05 ( 1000 993 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU05 ( 999 993 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU05 ( 998 993 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU05 ( 997 993 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU05 ( 996 993 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU05 ( 995 993 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU05 ( 994 993 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU05 ( 992 993 ) COMPLEX( 100.n, 0.)
R_D52132LOADxxU05 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U06CCM 
R_D52101xxU06 ( 1027 1059 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU06 ( 1058 1027 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU06 ( 1057 1027 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU06 ( 1056 1027 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU06 ( 1055 1027 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU06 ( 1054 1027 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxU06 ( 1053 1027 ) COMPLEX( 100.n, 0.)
R_D52107xxU06 ( 1052 1027 ) COMPLEX( 100.n, 0.)
R_D52109xxU06 ( 1051 1027 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU06 ( 1050 1027 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU06 ( 1049 1027 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU06 ( 1048 1027 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU06 ( 1047 1027 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU06 ( 1046 1027 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU06 ( 1045 1027 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxU06 ( 584 1027 ) COMPLEX( 100.n, 0.)
R_D52115xxU06 ( 1043 1027 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU06 ( 1027 1042 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU06 ( 1041 1027 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU06 ( 1040 1027 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU06 ( 1039 1027 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU06 ( 1038 1027 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU06 ( 1037 1027 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxU06 ( 1036 1027 ) COMPLEX( 100.n, 0.)
R_D52124xxU06 ( 1035 1027 ) COMPLEX( 100.n, 0.)
R_D52125xxU06 ( 1034 1027 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU06 ( 1033 1027 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU06 ( 1032 1027 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU06 ( 1031 1027 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU06 ( 1030 1027 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU06 ( 1029 1027 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU06 ( 1028 1027 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU06 ( 1026 1027 ) COMPLEX( 100.n, 0.)
R_D52132LOADxxU06 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*-------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U07CCM 
R_D52101xxU07 ( 1061 1093 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU07 ( 1092 1061 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU07 ( 1091 1061 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU07 ( 1090 1061 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU07 ( 1089 1061 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU07 ( 1088 1061 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxU07 ( 1087 1061 ) COMPLEX( 100.n, 0.)
R_D52107xxU07 ( 1086 1061 ) COMPLEX( 100.n, 0.)
R_D52109xxU07 ( 1085 1061 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU07 ( 1084 1061 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU07 ( 1083 1061 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU07 ( 1082 1061 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU07 ( 1081 1061 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU07 ( 1080 1061 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU07 ( 1079 1061 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxU07 ( 588 1061 ) COMPLEX( 100.n, 0.)
R_D52115xxU07 ( 1077 1061 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU07 ( 1061 1076 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU07 ( 1075 1061 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU07 ( 1074 1061 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU07 ( 1073 1061 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU07 ( 1072 1061 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU07 ( 1071 1061 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxU07 ( 1070 1061 ) COMPLEX( 100.n, 0.)
R_D52124xxU07 ( 1069 1061 ) COMPLEX( 100.n, 0.)
R_D52125xxU07 ( 1068 1061 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU07 ( 1067 1061 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU07 ( 1066 1061 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU07 ( 1065 1061 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU07 ( 1064 1061 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU07 ( 1063 1061 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU07 ( 1062 1061 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU07 ( 1060 1061 ) COMPLEX( 100.n, 0.)
R_D52132LOADxxU07 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*----------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA U08CCM 
R_D52101xxU08 ( 1095 1127 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxU08 ( 1126 1095 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxU08 ( 1125 1095 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxU08 ( 1124 1095 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxU08 ( 1123 1095 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxU08 ( 1122 1095 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxU08 ( 1121 1095 ) COMPLEX( 100.n, 0.)
R_D52107xxU08 ( 1120 1095 ) COMPLEX( 100.n, 0.)
R_D52109xxU08 ( 1119 1095 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxU08 ( 1118 1095 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxU08 ( 1117 1095 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxU08 ( 1116 1095 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxU08 ( 1115 1095 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxU08 ( 1114 1095 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxU08 ( 1113 1095 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52ExxU08 ( 587 1095 ) COMPLEX( 100.n, 0.)
R_D52115xxU08 ( 1111 1095 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52118xxU08 ( 1095 1110 ) COMPLEX( 100.n, 0.)
R_D52118LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52119xxU08 ( 1109 1095 ) COMPLEX( 100.n, 0.)
R_D52119LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52120xxU08 ( 1108 1095 ) COMPLEX( 100.n, 0.)
R_D52120LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52121xxU08 ( 1107 1095 ) COMPLEX( 100.n, 0.)
R_D52121LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52122xxU08 ( 1106 1095 ) COMPLEX( 100.n, 0.)
R_D52122LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52123xxU08 ( 1105 1095 ) COMPLEX( 100.n, 0.)
R_D52123LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52124LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52117xxU08 ( 1104 1095 ) COMPLEX( 100.n, 0.)
R_D52124xxU08 ( 1103 1095 ) COMPLEX( 100.n, 0.)
R_D52125xxU08 ( 1102 1095 ) COMPLEX( 100.n, 0.)
R_D52125LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52126xxU08 ( 1101 1095 ) COMPLEX( 100.n, 0.)
R_D52126LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52127xxU08 ( 1100 1095 ) COMPLEX( 100.n, 0.)
R_D52127LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52128xxU08 ( 1099 1095 ) COMPLEX( 100.n, 0.)
R_D52128LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52129xxU08 ( 1098 1095 ) COMPLEX( 100.n, 0.)
R_D52129LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52130xxU08 ( 1097 1095 ) COMPLEX( 100.n, 0.)
R_D52130LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52131xxU08 ( 1096 1095 ) COMPLEX( 100.n, 0.)
R_D52131LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52132xxU08 ( 1094 1095 ) COMPLEX( 100.n, 0.)
R_D52132LOADxxU08 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*---------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA CCME1 
R_D52E1xxCCME1 ( 583 1129 ) COMPLEX( 100.n, 0.)
R_D52E2xxCCME1 ( 597 1128 ) COMPLEX( 100.n, 0.)
R_D52206xxCCME1 ( 1142 1128 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxCCME1 ( 1141 1128 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxCCME1 ( 1140 1128 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxCCME1 ( 1139 1128 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxCCME1 ( 1138 1128 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxCCME1 ( 1137 1128 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxCCME1 ( 1136 1129 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxCCME1 ( 1135 1129 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxCCME1 ( 1134 1129 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxCCME1 ( 1133 1129 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxCCME1 ( 1132 1129 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxCCME1 ( 1131 1129 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxCCME1 ( 1130 1129 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52LxxCCME1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA CCME2 
R_D52E1xxCCME2 ( 572 1144 ) COMPLEX( 100.n, 0.)
R_D52E2xxCCME2 ( 565 1143 ) COMPLEX( 100.n, 0.)
R_D52206xxCCME2 ( 1157 1143 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxCCME2 ( 1156 1143 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxCCME2 ( 1155 1143 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxCCME2 ( 1154 1143 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxCCME2 ( 1153 1143 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxCCME2 ( 1152 1143 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxCCME2 ( 1151 1144 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxCCME2 ( 1150 1144 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxCCME2 ( 1149 1144 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxCCME2 ( 1148 1144 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxCCME2 ( 1147 1144 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxCCME2 ( 1146 1144 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxCCME2 ( 1145 1144 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52LxxCCME2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*---------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA CCMD1 
R_D52101xxCCMD1 ( 1180 1159 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52E1xxCCMD1 ( 454 1159 ) COMPLEX( 100.n, 0.)
R_D52209xxCCMD1 ( 1178 1169 ) COMPLEX( 100.n, 0.)
R_D52209LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52E2xxCCMD1 ( 595 1169 ) COMPLEX( 100.n, 0.)
R_D52208xxCCMD1 ( 1176 1169 ) COMPLEX( 100.n, 0.)
R_D52208LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207xxCCMD1 ( 1175 1169 ) COMPLEX( 100.n, 0.)
R_D52207LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxCCMD1 ( 1174 1169 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxCCMD1 ( 1173 1169 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxCCMD1 ( 1172 1169 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxCCMD1 ( 1171 1169 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxCCMD1 ( 1170 1169 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxCCMD1 ( 1168 1169 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxCCMD1 ( 1167 1159 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxCCMD1 ( 1166 1159 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxCCMD1 ( 1165 1159 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxCCMD1 ( 1164 1159 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxCCMD1 ( 1163 1159 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxCCMD1 ( 1162 1159 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxCCMD1 ( 1161 1159 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxCCMD1 ( 1160 1159 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxCCMD1 ( 1158 1159 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52LxxCCMD1 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*--------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA CCMD2 
R_D52101xxCCMD2 ( 1203 1182 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52E1xxCCMD2 ( 567 1182 ) COMPLEX( 100.n, 0.)
R_D52209xxCCMD2 ( 1201 1192 ) COMPLEX( 100.n, 0.)
R_D52209LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52E2xxCCMD2 ( 560 1192 ) COMPLEX( 100.n, 0.)
R_D52208xxCCMD2 ( 1199 1192 ) COMPLEX( 100.n, 0.)
R_D52208LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207xxCCMD2 ( 1198 1192 ) COMPLEX( 100.n, 0.)
R_D52207LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxCCMD2 ( 1197 1192 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxCCMD2 ( 1196 1192 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxCCMD2 ( 1195 1192 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxCCMD2 ( 1194 1192 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxCCMD2 ( 1193 1192 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxCCMD2 ( 1191 1192 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxCCMD2 ( 1190 1182 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxCCMD2 ( 1189 1182 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxCCMD2 ( 1188 1182 ) COMPLEX( 100.n, 0.)
R_D52108LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxCCMD2 ( 1187 1182 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxCCMD2 ( 1186 1182 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxCCMD2 ( 1185 1182 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxCCMD2 ( 1184 1182 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxCCMD2 ( 1183 1182 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxCCMD2 ( 1181 1182 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52LxxCCMD2 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSSE3 
R_D52E1xxQSSE3 ( 593 1206 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSSE3 ( 622 1209 ) COMPLEX( 100.n, 0.)
R_D52307xxQSSE3 ( 1218 1204 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSSE3 ( 1217 1204 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSSE3 ( 1216 1204 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSSE3 ( 1215 1204 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSSE3 ( 1214 1204 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSSE3 ( 1213 1204 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSSE3 ( 1212 1204 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSSE3 ( 1211 1209 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSSE3 ( 1210 1209 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSSE3 ( 1208 1209 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSSE3 ( 1207 1206 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSSE3 ( 1205 1206 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSSE3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L2xxQSSE3 ( 1204 1209 ) COMPLEX( 100.n, 0.)
*------------------------------------------------------------------------------------------------------------------------------------------------------------------ 
*Netlist: Auxiliares CA QSSE4 
R_D52E1xxQSSE4 ( 616 1221 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSSE4 ( 601 1225 ) COMPLEX( 100.n, 0.)
R_D52307xxQSSE4 ( 1234 1219 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSSE4 ( 1233 1219 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSSE4 ( 1232 1219 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSSE4 ( 1231 1219 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSSE4 ( 1230 1219 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSSE4 ( 1229 1219 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52301xxQSSE4 ( 1228 1219 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSSE4 ( 1227 1225 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSSE4 ( 1226 1225 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52201xxQSSE4 ( 1224 1225 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSSE4 ( 1223 1221 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSSE4 ( 1222 1221 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52101xxQSSE4 ( 1220 1221 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSSE4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L2xxQSSE4 ( 1219 1225 ) COMPLEX( 100.n, 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
*Netlist: Auxiliares CA QSG3 
R_D52101xxQSG3 ( 1241 1301 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSG3 ( 1300 1241 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSG3 ( 1299 1241 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSG3 ( 1298 1241 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSG3 ( 1297 1241 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxQSG3 ( 1296 1241 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxQSG3 ( 1295 1241 ) COMPLEX( 100.n, 0.)
R_D52110xxQSG3 ( 1294 1241 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52111xxQSG3 ( 1293 1241 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSG3 ( 1292 1241 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSG3 ( 1291 1241 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxQSG3 ( 1290 1241 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSG3 ( 1289 1241 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52116xxQSG3 ( 1287 1241 ) COMPLEX( 100.n, 0.)
R_D52116LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSG3 ( 1286 1241 ) COMPLEX( 100.n, 0.)
R_D52109LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L2xxQSG3 ( 1236 1267 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSG3 ( 618 1267 ) COMPLEX( 100.n, 0.)
R_D52E1xxQSG3 ( 592 1241 ) COMPLEX( 100.n, 0.)
R_D52201xxQSG3 ( 1267 1284 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSG3 ( 1283 1267 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSG3 ( 1282 1267 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQSG3 ( 1281 1267 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQSG3 ( 1280 1267 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQSG3 ( 1279 1267 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52208LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52208xxQSG3 ( 1278 1267 ) COMPLEX( 100.n, 0.)
R_D52210xxQSG3 ( 1277 1267 ) COMPLEX( 100.n, 0.)
R_D52210LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52211xxQSG3 ( 1276 1267 ) COMPLEX( 100.n, 0.)
R_D52211LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52212xxQSG3 ( 1275 1267 ) COMPLEX( 100.n, 0.)
R_D52212LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52213xxQSG3 ( 1274 1267 ) COMPLEX( 100.n, 0.)
R_D52213LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52214xxQSG3 ( 1273 1267 ) COMPLEX( 100.n, 0.)
R_D52214LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52215xxQSG3 ( 1272 1267 ) COMPLEX( 100.n, 0.)
R_D52215LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52216xxQSG3 ( 1271 1267 ) COMPLEX( 100.n, 0.)
R_D52216LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52209xxQSG3 ( 1270 1267 ) COMPLEX( 100.n, 0.)
R_D52209LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52326xxQSG3 ( 1269 1236 ) COMPLEX( 100.n, 0.)
R_D52326LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52327xxQSG3 ( 1268 1236 ) COMPLEX( 100.n, 0.)
R_D52327LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207xxQSG3 ( 1266 1267 ) COMPLEX( 100.n, 0.)
R_D52301xxQSG3 ( 1236 1264 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSG3 ( 1263 1236 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSG3 ( 1262 1236 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSG3 ( 1261 1236 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSG3 ( 1260 1236 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSG3 ( 1259 1236 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52308LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52308xxQSG3 ( 1258 1236 ) COMPLEX( 100.n, 0.)
R_D52311xxQSG3 ( 1257 1236 ) COMPLEX( 100.n, 0.)
R_D52311LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52312xxQSG3 ( 1256 1236 ) COMPLEX( 100.n, 0.)
R_D52312LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52313xxQSG3 ( 1255 1236 ) COMPLEX( 100.n, 0.)
R_D52313LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52314xxQSG3 ( 1254 1236 ) COMPLEX( 100.n, 0.)
R_D52314LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52315xxQSG3 ( 1253 1236 ) COMPLEX( 100.n, 0.)
R_D52315LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52316xxQSG3 ( 1252 1236 ) COMPLEX( 100.n, 0.)
R_D52316LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52317xxQSG3 ( 1251 1236 ) COMPLEX( 100.n, 0.)
R_D52317LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52310xxQSG3 ( 1250 1236 ) COMPLEX( 100.n, 0.)
R_D52310LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52318xxQSG3 ( 1249 1236 ) COMPLEX( 100.n, 0.)
R_D52318LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319xxQSG3 ( 1248 1236 ) COMPLEX( 100.n, 0.)
R_D52319LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309xxQSG3 ( 1247 1236 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52307xxQSG3 ( 1246 1236 ) COMPLEX( 100.n, 0.)
R_D52320xxQSG3 ( 1236 1245 ) COMPLEX( 100.n, 0.)
R_D52320LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52321xxQSG3 ( 1244 1236 ) COMPLEX( 100.n, 0.)
R_D52321LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52325xxQSG3 ( 1243 1236 ) COMPLEX( 100.n, 0.)
R_D52325LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52324xxQSG3 ( 1242 1236 ) COMPLEX( 100.n, 0.)
R_D52324LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSG3 ( 1240 1241 ) COMPLEX( 100.n, 0.)
R_D52322xxQSG3 ( 1238 1236 ) COMPLEX( 100.n, 0.)
R_D52322LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52323xxQSG3 ( 1237 1236 ) COMPLEX( 100.n, 0.)
R_D52323LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52328xxQSG3 ( 1235 1236 ) COMPLEX( 100.n, 0.)
R_D52328LOADxxQSG3 ( 0 0 ) COMPLEX( 1.E+12, 0.)
*----------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA QSG4 
R_D52101xxQSG4 ( 1346 1361 ) COMPLEX( 100.n, 0.)
R_D52101LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52102xxQSG4 ( 1360 1346 ) COMPLEX( 100.n, 0.)
R_D52102LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52103xxQSG4 ( 1359 1346 ) COMPLEX( 100.n, 0.)
R_D52103LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52104xxQSG4 ( 1358 1346 ) COMPLEX( 100.n, 0.)
R_D52104LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52105xxQSG4 ( 1357 1346 ) COMPLEX( 100.n, 0.)
R_D52105LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52107xxQSG4 ( 1356 1346 ) COMPLEX( 100.n, 0.)
R_D52107LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52108xxQSG4 ( 1355 1346 ) COMPLEX( 100.n, 0.)
R_D52111xxQSG4 ( 1354 1346 ) COMPLEX( 100.n, 0.)
R_D52111LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52112xxQSG4 ( 1353 1346 ) COMPLEX( 100.n, 0.)
R_D52112LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52113xxQSG4 ( 1352 1346 ) COMPLEX( 100.n, 0.)
R_D52113LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52114xxQSG4 ( 1351 1346 ) COMPLEX( 100.n, 0.)
R_D52114LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52115xxQSG4 ( 1350 1346 ) COMPLEX( 100.n, 0.)
R_D52115LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52L1xxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52110xxQSG4 ( 1348 1346 ) COMPLEX( 100.n, 0.)
R_D52110LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52109xxQSG4 ( 1347 1346 ) COMPLEX( 100.n, 0.)
R_D52106LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52106xxQSG4 ( 1345 1346 ) COMPLEX( 100.n, 0.)
R_D52L2xxQSG4 ( 1303 1327 ) COMPLEX( 100.n, 0.)
R_D52E2xxQSG4 ( 598 1327 ) COMPLEX( 100.n, 0.)
R_D52E1xxQSG4 ( 614 1346 ) COMPLEX( 100.n, 0.)
R_D52201xxQSG4 ( 1327 1342 ) COMPLEX( 100.n, 0.)
R_D52201LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52202xxQSG4 ( 1341 1327 ) COMPLEX( 100.n, 0.)
R_D52202LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52203xxQSG4 ( 1340 1327 ) COMPLEX( 100.n, 0.)
R_D52203LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52204xxQSG4 ( 1339 1327 ) COMPLEX( 100.n, 0.)
R_D52204LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52205xxQSG4 ( 1338 1327 ) COMPLEX( 100.n, 0.)
R_D52205LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52206xxQSG4 ( 1337 1327 ) COMPLEX( 100.n, 0.)
R_D52206LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52208LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52208xxQSG4 ( 1336 1327 ) COMPLEX( 100.n, 0.)
R_D52211xxQSG4 ( 1335 1327 ) COMPLEX( 100.n, 0.)
R_D52211LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52212xxQSG4 ( 1334 1327 ) COMPLEX( 100.n, 0.)
R_D52212LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52213xxQSG4 ( 1333 1327 ) COMPLEX( 100.n, 0.)
R_D52213LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52214xxQSG4 ( 1332 1327 ) COMPLEX( 100.n, 0.)
R_D52214LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52215xxQSG4 ( 1331 1327 ) COMPLEX( 100.n, 0.)
R_D52215LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52216xxQSG4 ( 1330 1327 ) COMPLEX( 100.n, 0.)
R_D52216LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52210xxQSG4 ( 1329 1327 ) COMPLEX( 100.n, 0.)
R_D52210LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52209LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52209xxQSG4 ( 1328 1327 ) COMPLEX( 100.n, 0.)
R_D52207LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52207xxQSG4 ( 1326 1327 ) COMPLEX( 100.n, 0.)
R_D52301xxQSG4 ( 1303 1324 ) COMPLEX( 100.n, 0.)
R_D52301LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52302xxQSG4 ( 1323 1303 ) COMPLEX( 100.n, 0.)
R_D52302LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52303xxQSG4 ( 1322 1303 ) COMPLEX( 100.n, 0.)
R_D52303LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52304xxQSG4 ( 1321 1303 ) COMPLEX( 100.n, 0.)
R_D52304LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52305xxQSG4 ( 1320 1303 ) COMPLEX( 100.n, 0.)
R_D52305LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52306xxQSG4 ( 1319 1303 ) COMPLEX( 100.n, 0.)
R_D52306LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52308LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52308xxQSG4 ( 1318 1303 ) COMPLEX( 100.n, 0.)
R_D52311xxQSG4 ( 1317 1303 ) COMPLEX( 100.n, 0.)
R_D52311LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52312xxQSG4 ( 1316 1303 ) COMPLEX( 100.n, 0.)
R_D52312LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52313xxQSG4 ( 1315 1303 ) COMPLEX( 100.n, 0.)
R_D52313LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52314xxQSG4 ( 1314 1303 ) COMPLEX( 100.n, 0.)
R_D52314LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52315xxQSG4 ( 1313 1303 ) COMPLEX( 100.n, 0.)
R_D52315LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52316xxQSG4 ( 1312 1303 ) COMPLEX( 100.n, 0.)
R_D52316LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52317xxQSG4 ( 1311 1303 ) COMPLEX( 100.n, 0.)
R_D52317LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52310xxQSG4 ( 1310 1303 ) COMPLEX( 100.n, 0.)
R_D52310LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52318xxQSG4 ( 1309 1303 ) COMPLEX( 100.n, 0.)
R_D52318LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52319xxQSG4 ( 1308 1303 ) COMPLEX( 100.n, 0.)
R_D52319LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52309xxQSG4 ( 1307 1303 ) COMPLEX( 100.n, 0.)
R_D52307LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52307xxQSG4 ( 1306 1303 ) COMPLEX( 100.n, 0.)
R_D52320xxQSG4 ( 1303 1305 ) COMPLEX( 100.n, 0.)
R_D52320LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52321xxQSG4 ( 1304 1303 ) COMPLEX( 100.n, 0.)
R_D52321LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52322LOADxxQSG4 ( 0 0 ) COMPLEX( 1.E+12, 0.)
R_D52322xxQSG4 ( 1302 1303 ) COMPLEX( 100.n, 0.)
*-------------------------------------------------------------------------------------------------------------------------------------------------------------- 
* Netlist: Auxiliares CA U09CCM 
.end